Require Import List.

Require Import Logic.Class.Eq.

Require Import Logic.Func.Permute.
Require Import Logic.Func.Identity.
Require Import Logic.Func.Injective.
Require Import Logic.Func.Composition.

Require Import Logic.List.In.
Require Import Logic.List.Remove.
Require Import Logic.List.Append.
Require Import Logic.List.InjectiveOn.

Require Import Logic.Lam.Free.
Require Import Logic.Lam.Valid.
Require Import Logic.Lam.Syntax.
Require Import Logic.Lam.Functor.
Require Import Logic.Lam.Variable.
Require Import Logic.Lam.Congruence.
Require Import Logic.Lam.Admissible.

(* Generator of alpha-equivalence.                                              *)
(* We wish to formally define alpha-equivalence as the smallest congruence      *)
(* contaning all ordered pairs below. Note that we are using the permutation    *)
(* y <:> x rather than the substitution (y // x) and we allow the variable y    *)
(* to be a variable of t1 as long as it is not free. This seemingly unusual     *)
(* choice is to make sure we obtain a definition of alpha-equivalence which     *)
(* works equally well for a finite or infinite variable type v. Otherwise, we   *)
(* would obtain a congruence which is strictly stronger than alpha-equivalence  *)
(* when v is finite. See the StrongAlpha module for details.                    *)
Inductive Alpha0 (v:Type) (e:Eq v) : T v -> T v -> Prop :=
| mkAlpha0: forall (x y:v) (t1:T v), 
    x <> y       -> 
    ~ y :: Fr t1 ->
    Alpha0 v e (Lam x t1) (Lam y (fmap (y <:> x) t1)) 
.

Arguments Alpha0 {v} {e}.
Arguments mkAlpha0 {v} {e}.

(* The alpha-equivalence relation is the congruence generated by Alph0.         *)
Definition Alpha (v:Type) (e:Eq v) : T v -> T v -> Prop := 
    Cong (@Alpha0 v e).

Arguments Alpha {v} {e}.

Notation "t ~ s" := (Alpha t s)
    (at level 60, no associativity) : Lam_Alpha_scope.

Open Scope Lam_Alpha_scope.

(* Admissible substitutions do not change alpha-equivalence classes.            *)
Lemma Alpha_admissible : forall (v:Type) (e:Eq v) (t:T v) (f:v -> v),
  admissible f t -> t ~ fmap f t.
Proof.
  intros v e.
  induction t as [x|t1 IH1 t2 IH2|x t1 IH1]; 
  intros f [H1 H2]; simpl; simpl in H2.

  (* case t = Var x *)
  - assert (f x = x) as E1. { apply H2. left. reflexivity. }
    rewrite E1. apply Cong_reflexive.

  (* case t = App t1 t2 *)
  - rewrite valid_app in H1; destruct H1 as [H1 H3].

    assert (t1 ~ fmap f t1) as E1.
      { apply IH1. unfold admissible. split.
        { assumption. }
        { intros x H4. apply H2, app_charac. left. assumption. }}

    assert (t2 ~ fmap f t2) as E2.
      { apply IH2. unfold admissible. split.
        { assumption. }
        { intros x H4. apply H2, app_charac. right. assumption. }}

    apply CongApp; assumption. 

  (* case t = Lam x t1 *)
  - rewrite valid_lam in H1. destruct H1 as [H3 H4].
    destruct (eqDec (f x) x) as [H5|H5].

    + (* f x = x *)
      assert (t1 ~ fmap f t1) as E1.
        { apply IH1. unfold admissible. split.
          { assumption. }
          { intros y H6.
            assert (f y = y) as E1.
              { destruct (eqDec x y) as [H7|H7].
                { (* x = y  *)
                  rewrite <- H7. assumption. }
                { (* x <> y *)
                  apply H2, remove_charac. split; assumption. }}
           assumption. }} 
      rewrite H5. apply CongLam. assumption.
      
    + (* f x <> x *)
      remember (f x) as y eqn:H6.

      assert (Lam x t1 ~ Lam y (fmap f t1)) as E.
        { remember ((y <:> x) ; f) as g eqn:H7.
          remember (fmap g t1) as s1 eqn:H8. 

          assert (f = (y <:> x) ; g) as E1.
            { rewrite H7. rewrite comp_assoc, permute_involution.
              symmetry. apply comp_id_left. }

          assert (fmap f t1 = fmap (y <:> x) s1) as E2.
            { rewrite H8, <- fmap_comp', <- E1. reflexivity. }

          rewrite E2.

          assert (Lam x t1 ~ Lam y (fmap (y <:> x) s1)) as E3.
            { assert (admissible g t1) as E8. 
                { unfold admissible. split.
                   { rewrite H7. rewrite <- valid_compose. split.
                    { apply H3. (* why is the assumption tactic failing here *) }
                    { apply valid_inj, injective_injective_on. 
                      apply permute_injective. }}
                { intros u H10. destruct (eqDec u x) as [H11|H11].
                    { subst. unfold comp. apply permute_app_left. }
                    { rewrite H7. unfold comp. 
                      assert (f u = u) as H12.
                        { apply H2. apply remove_charac. split.
                          { assumption. }
                          { intros H12. apply H11. symmetry.  assumption. }}
                      rewrite H12. apply permute_app_diff. 
                        { intros H13. apply H4 with u. 
                          { simpl. apply remove_charac. split.
                            { assumption. }
                            { intros H14. apply H11. symmetry. assumption. }}
                          { rewrite H12. symmetry. assumption. }}
                        { assumption. }}}}

              assert (~ y :: Fr s1) as E4.
                { rewrite H8. intros H9. apply (free_fmap v v e) in H9.
                  apply in_map_iff in H9. destruct H9 as [u [H9 H10]].
                  unfold admissible in E8. destruct E8 as [H11 H12]. 
        
                  assert (g u = u) as H13. { apply H12. assumption. }

                  assert (y :: Fr t1) as H14. { rewrite <- H9, H13. assumption. }
              
                  assert (y :: Fr (Lam x t1)) as H15.
                    { simpl. apply remove_charac. split.
                      { assumption. }
                      { intros H16. apply H5. symmetry. assumption. }} 

                  assert (f y = y) as H17. { apply H2. assumption. }

                  assert (f x <> f y) as H18. 
                    { rewrite <- H6. apply H4. assumption. }

                  assert (f x <> y) as H19. { rewrite <- H17. assumption. }
  
                  apply H19. symmetry. assumption. }

              assert (Lam x s1 ~ Lam y (fmap (y <:> x) s1)) as E5.
                { constructor. constructor.
                  { intros H9. apply H5. symmetry. assumption. }
                  { assumption. }}

              assert (Lam x t1 ~ Lam x s1) as E6.
                { assert (t1 ~ s1) as E7. { rewrite H8. apply IH1. apply E8. }
                  apply Cong_congruent, E7. }

              apply Cong_transitive with (Lam x s1); assumption. }
          apply E3. }
      apply E.
Qed.
