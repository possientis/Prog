Require Import List.

Require Import Logic.Class.Eq.

Require Import Logic.Rel.R.
Require Import Logic.Rel.Include.

Require Import Logic.Func.Permute.
Require Import Logic.Func.Identity.
Require Import Logic.Func.Injective.
Require Import Logic.Func.Composition.

Require Import Logic.List.In.
Require Import Logic.List.Remove.
Require Import Logic.List.Append.
Require Import Logic.List.Coincide.
Require Import Logic.List.InjectiveOn.

Require Import Logic.Lam.Free.
Require Import Logic.Lam.Valid.
Require Import Logic.Lam.Syntax.
Require Import Logic.Lam.Functor.
Require Import Logic.Lam.Variable.
Require Import Logic.Lam.Congruence.
Require Import Logic.Lam.Subformula.
Require Import Logic.Lam.Admissible.

Declare Scope Lam_Alpha_scope.

(* Generator of alpha-equivalence.                                              *)
(* We wish to formally define alpha-equivalence as the smallest congruence      *)
(* contaning all ordered pairs below. Note that we are using the permutation    *)
(* y <:> x rather than the substitution (y // x) and we allow the variable y    *)
(* to be a variable of t1 as long as it is not free. This seemingly unusual     *)
(* choice is to make sure we obtain a definition of alpha-equivalence which     *)
(* works equally well for a finite or infinite variable type v. Otherwise, we   *)
(* would obtain a congruence which is strictly stronger than alpha-equivalence  *)
(* when v is finite. See the StrongAlpha module for details.                    *)
Inductive Alpha0 (v:Type) (e:Eq v) : T v -> T v -> Prop :=
| mkAlpha0: forall (x y:v) (t1:T v), 
    x <> y       -> 
    ~ y :: Fr t1 ->
    Alpha0 v e (Lam x t1) (Lam y (fmap (y <:> x) t1)) 
.

Arguments Alpha0 {v} {e}.
Arguments mkAlpha0 {v} {e}.

(* The alpha-equivalence relation is the congruence generated by Alph0.         *)
Definition Alpha (v:Type) (e:Eq v) : T v -> T v -> Prop := 
    Cong (@Alpha0 v e).

Arguments Alpha {v} {e}.

Notation "t ~ s" := (Alpha t s)
    (at level 60, no associativity) : Lam_Alpha_scope.

Open Scope Lam_Alpha_scope.

(* Admissible substitutions do not change alpha-equivalence classes.            *)
Lemma Alpha_admissible : forall (v:Type) (e:Eq v) (t:T v) (f:v -> v),
  admissible f t -> t ~ fmap f t.
Proof.
  (* Let v be a Type with decidable equality e  *)
  intros v e.

  (* We prove the lemma with an induction argument on t *)
  induction t as [x|t1 IH1 t2 IH2|x t1 IH1]; 

  (* In each case we assume f:v -> v is valid for t with f u = u for u :: Fr t  *)
  intros f H1.

  (* case t = Var x *)
  - assert (Var x ~ Var (f x)) as A. 2: apply A.

    assert (f x = x) as A1. 
    { apply admissible_free with (Var x).
      - apply H1.
      - left. reflexivity.
    }

    rewrite A1.

    apply Cong_reflexive.

  (* case t = App t1 t2 *)
  - assert (App t1 t2 ~ App (fmap f t1) (fmap f t2)) as A. 2: apply A. 

    (* Note that f being admissible for App t1 t2  ... *)
    apply admissible_app in H1. destruct H1 as [H1 H2].
    
    (* ... it is admissible for t1 ... *)
    assert (admissible f t1) as A. apply H1. clear A.

    (* ... and it is admissible for t2 *)
    assert (admissible f t2)as A. apply H2. clear A.


    (* We argue that alpha-equivalence is a congruence  *)
    apply CongApp.

    (* So we need to prove that t1 ~ fmap f t1  *)
    + assert (t1 ~ fmap f t1) as A. 2: apply A. 

      (* This follows from the induction hypothesis ... *)
      apply IH1. 

      (* ... provided we show that f is admissible for t1 *)
      assert (admissible f t1) as A. 2: apply A.
 
      (* ... which we know is true  *) 
      apply H1.

    (* We need to prove similarly that t2 ~ fmap f t2  *)
    + assert (t2 ~ fmap f t2) as A. 2: apply A.

      (* This follows from the induction hypothesis ... *)
      apply IH2.

      (* ... provided we show that f is admissible for t2 *)
      assert (admissible f t2) as A. 2: apply A.

      (* ... which we know is true *)
      apply H2.

  (* case p = Lam x t1 *)
  - assert (Lam x t1 ~ Lam (f x) (fmap f t1)) as A. 2: apply A. 

    (* Note that f being admissible for Lam x t1 ... *)
    destruct H1 as [H1 H3]. apply valid_lam in H1. destruct H1 as [H1 H2].

    (* ... it is valid for t1 ... *)
    assert (valid f t1) as A. apply H1. clear A.

    (* ... we have f x <> f y for any y free in Lam x t1  ... *)
    assert (forall (y:v), y :: Fr (Lam x t1)->f x <> f y) as A. apply H2. clear A.

    (* ... and we have f y = y for any y free in Lam x t1 *)
    assert (forall (y:v), y :: Fr (Lam x t1) -> f y = y) as A. apply H3. clear A.
 
    (* We carry out the proof by distinguishing two cases *)
    destruct (eqDec (f x) x) as [H4|H4].

    + (* First we assume that f x = x *)

      (* Given that f x = x *)
      rewrite H4.

      (* We need to show that Lam x t1 ~ Lam x (fmap f t1)  *)
      assert (Lam x t1 ~ Lam x (fmap f t1)) as A. 2: apply A.

      (* Alpha-equivalence being a congruence ... *)
      apply CongLam.

      (* ... we simply need to show that t1 ~ fmap f t1 *)
      assert (t1 ~ fmap f t1) as A. 2: apply A.

      (* This follows from the induction hypothesis ... *)
      apply IH1.

      (* ... provided we show that f is admissible for t1 *)
      assert (admissible f t1) as A. 2: apply A.

      (* Given the definition of an admissible mapping ... *)
      unfold admissible. split.

      (* ... we need to show that f is valid for t1 ... *)
      * assert (valid f t1) as A. 2: apply A.

        (* ... which is true as we have noted *)
        apply H1.

      (* ... and that free variables of t1 are invariant by f *)
      * assert (forall (u:v), u :: Fr t1 -> f u = u) as A. 2: apply A.

        (* So let u with u :: Fr t1 *)
        intros u H5. 
      
        (* We need to show that f u = u ... *) 
        assert (f u = u) as A. 2: apply A.

        (* We shall distinguish two cases *)
        destruct (eqDec x u) as [H6|H6].

        (* First we assume that x = u *)
        { rewrite <- H6.

          (* Then we need to show that f x = x ...  *)
          assert (f x = x) as A. 2: apply A.

          (* ... which we have assumed is true. *)
          apply H4.
        }

        (* Next we assume that x <> u *)
        { 
          (* Then f u = u follows from H3 ...*)
          apply H3.

          (* ... provided we show that u is free in Lam x t1  *) 
          assert (u :: Fr (Lam x t1)) as A. 2: apply A.
           
          simpl. apply remove_charac. split; assumption.
        }

    + (* Then we assume that f x <> x *)

      (* Define y *)
      remember (f x) as y eqn:E1.

      (* Define g *)
      remember ((y <:> x) ; f) as g eqn:E2.

      (* Define s1  *)
      remember (fmap g t1) as s1 eqn:E3. 

      (* So we need to show:  *)
      assert (Lam x t1 ~ Lam y (fmap f t1)) as A. 2: apply A.

      (* We claim that: *)
      assert (f = (y <:> x) ; g) as A1.
      { rewrite E2, comp_assoc, permute_involution. 
        symmetry. apply comp_id_left. 
      }
    
      (* And furthermore: *) 
      assert (fmap f t1 = fmap (y <:> x) s1) as A2.
      { rewrite E3, <- fmap_comp', <- A1. clear A1. reflexivity. 
      }

      (* We also claim that g is admissible for t1  *)
      assert (admissible g t1) as A3.
      { (* Given the definition of an admissible mapping ... *)
        unfold admissible. split.

        (* ... need need to show that g is valid for t1 *)
        - assert (valid g t1) as A. 2: apply A.

          (* Since g = (y <:> x) ; f  ... *)
          rewrite E2. 

          (* ... we need to show: *)
          assert (valid ((y <:> x) ; f) t1) as A. 2: apply A.

          (* and consequently ... *)
          rewrite <- valid_compose. split.

          (* ... we need to show that f is valid for t1 ... *)
          +  assert (valid f t1) as A. 2: apply A.
            
             (* ... we which know is true *)
             apply H1.

          (* ... and we need to show that (y <:> x) is valid for fmap f t1 ...*)
          + assert (valid (y <:> x) (fmap f t1)) as A. 2: apply A.

            (* ... which follows from the injectivity of pernutations *)
            apply valid_inj, injective_injective_on, permute_injective.

        (* ... and show that free variables of t1 are invariant by g  *)
        - assert (forall (u:v), u :: Fr t1 -> g u = u) as A. 2: apply A.

          (* so let u with u :: Fr t1 *)
          intros u H5. 

          (* We need to show that g u = u *)
          assert (g u = u) as A. 2: apply A.

          (* Given that g = (y <:> x) ... *)
          rewrite E2. unfold comp.

          (* ... amounts to showing that: *)
          assert ((y <:> x) (f u) = u) as A. 2: apply A.

          (* We shall distinguish two cases *)
          destruct (eqDec u x) as [H6|H6].

          * (* We first assume that u = x *)

            (* Given that u = x and y = f x ... *)
            rewrite H6, E1.

            (* ... we need to show that:  *)
            assert ((f x <:> x) (f x) = x) as A. 2: apply A.

            (* This is an immediate property of the permutation mapping *)
            apply permute_app_left.

          * (* We then assume that u <> x *)

            (* We claim that f u = u *)
            assert (f u = u) as A4.
            { (* This follows from H3 ... *)  
              apply H3. 

              (* ... provided we show that u is free in Lam x t1  *)
              assert (u :: Fr (Lam x t1)) as A. 2: apply A.

              simpl. apply remove_charac. split.

              (* So we need to show that u is free in t1 ...  *)
              - assert (u :: Fr t1) as A. 2: apply A.
                    
                apply H5.
              
              (* ... and that x <> u  *)
              - assert (x <> u) as A. 2: apply A.

                apply not_eq_sym, H6. 
            }

            (* So given that f u = u ... *)
            rewrite A4.

            (* we need to show that:  *)
            assert ((y <:> x) u = u) as A. 2: apply A.

            (* Hence, it is sufficient to prove... *)
            apply permute_app_diff.

            (* ... that u <> y  *)
            { assert (u <> y) as A. 2: apply A.

              (* So suppose that u = y  *)
              intros H7.

              (* Then we obtain a contradiction by showing f u <> u *)
              assert (f u <> u) as A. 2: contradiction.

              (* Given that u = y ... *)
              apply not_eq_sym. rewrite H7 at 1.

              (* ... we need to show that y <> f u  *)
              assert (y <> f u) as A. 2: apply A. 

              (* This follows from H2 ... *)
              apply H2.

              (* ... provided we show that u is free in Lam x t1 *)
              assert (u :: Fr (Lam x t1)) as A. 2: apply A.
         
              simpl. apply remove_charac. split.

              (* So we need to show that u is free in t1 ...  *)
              - assert (u :: Fr t1) as A. 2: apply A.
                  
                apply H5.

              (* ... and that x <> u  *)
              - assert (x <> u) as A. 2: apply A. 
                
                apply not_eq_sym, H6. 
            }

            (* ... and u <> x  *)
            { assert (u <> x) as A. 2: apply A.
                  
              apply H6.
            }
      (* This completes the proof of the admissibility of g for t1  *)
      } 

      (* So we now need to show:  *)
      assert (Lam x t1 ~ Lam y (fmap f t1)) as A. 2: apply A.

      (* Given that fmap f t1 = fmap (y <:> x) s1 ... *)
      rewrite A2. clear A2.

      (* ... we need to show that:  *)
      assert (Lam x t1 ~ Lam y (fmap (y <:> x) s1)) as A. 2: apply A.

      (* Alpha-equivalence being a transitive relation ...  *)
      apply Cong_transitive with (Lam x s1).

      (* ... it is sufficient to show firstly that: *) 
      * assert (Lam x t1 ~ Lam x s1) as A. 2: apply A.

        (* Alpha-equivalence being a congruence ... *)
        apply Cong_congruent.

        (* ... it is sufficient to show that t1 ~ s1 *)
        assert (t1 ~ s1) as A. 2: apply A.

        (* Given that s1 = fmap g t1  *)
        rewrite E3.

        (* we need to show that t1 ~ fmap q t1 ... *)
        assert (t1 ~ fmap g t1) as A. 2: apply A.

        (* ... which follows from the induction hypothesis ... *)
        apply IH1.

        (* ... provided we show show that g is admissible for t1 ...  *)
        assert (admissible g t1) as A. 2: apply A.

        (* ... which we have already proven *)
        apply A3.

      (* ... and secondly that:  *)
      * assert (Lam x s1 ~ Lam y (fmap (y <:> x) s1)) as A. 2: apply A.

        (* We argue that the pair actually belongs to the generator Alpha0  *)
        constructor.

        (* So we need to show that: *)
        assert (Alpha0 (Lam x s1) (Lam y (fmap (y <:> x) s1))) as A. 2: apply A.

        (* This is true by definition ...  *)
        constructor.

        (* ... provided we show that x <> y ... *)
        { assert (x <> y) as A. 2: apply A. 
          
          (* ... which is true since with have assumed f x <> x *)
          apply not_eq_sym, H4.
        }

        (* ... and that y is not free in s1 *)
        { assert (~ y :: Fr s1) as A. 2: apply A. 

          (* Given that s1 = fmap g t1 ...  *)
          rewrite E3. 

          (* ... we need to show that y is not free in fmap g t1 *)
          assert (~ y :: Fr (fmap g t1)) as A. 2: apply A. 

          (* So suppose to the contrary that y is free in fmap g t1 *)
          intros H5. 

          (* We need to obtain a contradiction by showing y <> f x *)
          assert (y <> f x) as A. 2: contradiction.

          (* Since Fr (fmap g t1) <= map g (Fr t1), we have y :: map g (Fr t1)  *)
          apply (free_fmap v v e) in H5.

          (* So there exists u such that y = g u and u :: Fr t1 *)
          apply in_map_iff in H5. destruct H5 as [u [H5 H6]].

          (* Note that g is valid for t1 and g u = u for all u :: Fr t1  *)
          unfold admissible in A3. destruct A3 as [H7 H8]. 

          (* It follows that g u = u *)
          assert (g u = u) as A4. { apply H8, H6. }

          (* It follows that y = u  *)
          assert (y = u) as A5. { rewrite <- A4. symmetry. apply H5. }

          (* So y is free in t1 *)
          assert (y :: Fr t1) as A6. { rewrite A5. apply H6. }

          (* So y is free in Lam x t1 *)
          assert (y :: Fr (Lam x t1)) as A7.
          { simpl. apply remove_charac. split.

            - assert (y :: Fr t1) as A. 2:apply A. apply A6.

            - assert (x <> y) as A. 2:apply A. apply not_eq_sym, H4.             
          }
         
          (* Hence from H3  we have f y = y *)
          assert (f y = y) as A8. { apply H3, A7. }

          (* Given that f y = y and y = f x ... *)
          rewrite <- A8, <- E1. apply not_eq_sym.

          (* We therefore need to show that y <> f y ... *) 
          assert (y <> f y) as A. 2: apply A.

          (* ... which follows from H2 ... *)
          apply H2. 

          (* ... provided we show that y is free in Lam x t1 ...  *)
          assert (y :: Fr (Lam x t1)) as A. 2: apply A.

          (* ... which has already been  established  *)
          apply A7.

        (* Completes the proof that y is not free in q1 *) 
        } 
Qed.

(* This is a relation which is larger than Alpha0 but a lot simpler. As we      *)
(* shall see, it is also a generator of the alpha-equivalence congruence.       *)
Inductive Alpha1 (v:Type) (e:Eq v) : T v -> T v -> Prop :=
| mkAlpha1: forall (t:T v) (f:v -> v), admissible f t -> Alpha1 v e t (fmap f t)
.

Arguments Alpha1 {v} {e}.
Arguments mkAlpha1 {v} {e}.

(* Alpha-equivalence is also the congruence generated by Alpha1.                *)
Lemma Alpha_admissible_gen : forall (v:Type) (e:Eq v), Alpha = Cong Alpha1.
Proof.
  (* Let v be a Type with decidable equality e  *)
  intros v e.
  
  (* Define r  *)
  remember (Cong Alpha1) as r eqn:E1.

  (* We need to show that Alpha = r *)
  assert (Alpha = r) as A. 2: apply A.

  (* We do so with a double inclusion argument *)
  apply incl_anti.

  (* First we show that Alpha <= r  *)
  - assert (Alpha <= r) as A. 2: apply A.

    (* We argue that Alpha is the smallest congruence containing Alpha0 *)
    unfold Alpha. apply Cong_smallest.

    (* So we need to show that r is a congruence  *)
    + assert (congruence r) as A. 2: apply A.
        
      rewrite E1. apply Cong_congruence.

    (* And we need to show that r contains Alpha0 *)
    + assert (Alpha0 <= r) as A. 2: apply A.

      (* So let x y and t1 such that x <> y and ~ y :: Fr t1  *)
      apply incl_charac. intros t s H1. destruct H1 as [x y t1 H1 H2].

      (* Define t *)
      remember (Lam x t1) as t eqn:E2.

      (* Define s *)
      remember (Lam y (fmap (y <:> x) t1)) as s eqn:E3.

      (* Define f *)
      remember (y <:> x) as f eqn:E4.

      (* We need to show that (p,q) :: r  *)
      assert (r t s) as A. 2: apply A.

      (* i.e. that (p.q) belongs to the congruence generated by Alpha1  *)
      rewrite E1. 
        
      (* We argue that (p,q) actually belongs to the generator itself *)
      constructor.

      (* So we need to show that (t,s) belongs to Alpha1  *)
      assert (Alpha1 t s) as A. 2: apply A.

      (* However, s is in fact s = fmap f t *)
      assert (s = fmap f t) as A.
      { rewrite E2, E3. simpl.
        assert (f x = y) as A5. 2: rewrite A5; reflexivity.
        rewrite E4. apply permute_app_right.
      }

      (* So we need to show that (t, fmap f t) lies in Alpha1 *)
      rewrite A. clear A. 
          
      (* which is true by definition... *)
      constructor.  
 
      (* ... provided we show that f is admissible for t  *)
      assert (admissible f t) as A. 2: apply A.

      (* Given the definition of an admissible substitution *)
      unfold admissible. split. 

      (* First we need to show that f is valid for t *)
      * assert (valid f t) as A. 2: apply A.
            
        (* It is sufficient to show that f is injective on (var t) *)
        apply valid_inj.
            
        (* It is sufficient to show that f is injective *)
        apply injective_injective_on.

        (* So we now prove that f is injective *)
        assert (injective f) as A. 2: apply A. 
            
        (* However, f is the permutation mapping (y <:> x)  *) 
        rewrite E4. 
            
        (* it is therefore injective  *)
        apply permute_injective.
         

      (* And furthermore that free variables are invariant by f *)
      * assert (forall (u:v), u :: Fr t -> f u = u) as A. 2: apply A.

        (* So let u with u :: Fr t  *) 
        intros u H3.
            
        (* We need to show that f u = u *)
        assert (f u = u) as A. 2: apply A.

        (* Given that f is the permutation mapping (y <:> x) ...  *)
        rewrite E4.

        (* ... it is sufficient to show that u <> x and u <> y *)
        apply permute_app_diff. 

        (* First we show that u <> y  *)
        { assert (u <> y) as A. 2: apply A.

          (* Since u :: Fr t, we have u :: Fr t1  *)
          assert (u :: Fr t1) as A.
          { rewrite E2 in H3. simpl in H3.
            apply remove_charac in H3.
            destruct H3 as [H3 H4]. assumption. 
          }
                
          (* So if we assume that u = y ... *)
          intros H4. 

          (* ... we obtain y :: Fr t1 which is a contradiction  *)
          rewrite H4 in A. contradiction. 
        }

        (* We now show that u <> x  *)
         { assert (u <> x) as A. 2: apply A.

          (* This is the case since u is free in p = All x p1 *)
          rewrite E2 in H3. simpl in H3. 
          apply remove_charac in H3.
          destruct H3 as [H3 H4]. apply not_eq_sym.
          assumption.

        } 
 
  (* We now show that r <= Alpha  *)
  - assert (r <= Alpha) as A. 2: apply A.

    (* We argue that r is the smallest congruence containing Alpha1 *)
    rewrite E1. apply Cong_smallest.

    (* So we need to show that Alpha is a congruence  *)
    + assert (congruence Alpha) as A. 2: apply A.
      
      unfold Alpha. apply Cong_congruence.
 
    (* And we need to show that Alpha contains Alpha1 *)
    + assert (Alpha1 <= Alpha) as A. 2: apply A.
      
      (* So let t and f : v -> v such that f is admissible for t  *) 
      apply incl_charac. intros t s H5. destruct H5 as [t f H5].

      (* We need to show that t is alpha-equivalent to fmap f t  *)
      assert (t ~ fmap f t) as A. 2: apply A. 

      (* This is the case, provided f is admissible for t ... *)
      apply Alpha_admissible. 
      
      (* ... which is true by assumption *)
      apply H5.
Qed.

(* Two alpha-equivalent formulas have the same free variables.                  *)
Lemma Alpha_free : forall (v:Type) (e:Eq v) (t s:T v), 
    t ~ s -> Fr t = Fr s.
Proof.
  (* Let v be a Type with decidable equality e  *)
  intros v e.  

  (* Define r to be the relation 'Fr t = Fr s' *)
  remember (fun (t s:T v) => Fr t = Fr s) as r eqn:E1.

  apply incl_charac. rewrite <- E1.

  (* We need to show that Alpha <= r  *)
  assert (Alpha <= r) as A. 2: apply A.

  (* We argue that Alpha is the smallest congruence containing Alpha1 *)
  rewrite Alpha_admissible_gen. apply Cong_smallest.

  (* So we need to show that r is a congruence ... *)
  - assert (congruence r) as A. 2: apply A.

    rewrite E1. apply free_congruence.

  (* ... and we need to show that r contains Alpha1 *)
  - assert (Alpha1 <= r) as A. 2: apply A.

    (* So let t be a formula and f:v -> v admissible for t *)
    apply incl_charac. intros t s H1. destruct H1 as [t f H1].
    
    (* We need to show that (t, fmap f t) lies in r *)
    assert (r t (fmap f t)) as A. 2: apply A.

    (* Given the way we have defined r ...  *)
    rewrite E1.

    (* ,,, we need to show that t and fmap f t have the same free variables *)
    assert (Fr t = Fr (fmap f t)) as A. 2: apply A.

    (* By transitivity ...  *)
    apply eq_trans with (map f (Fr t)).

    (* ... it is sufiicient to show firstly that Fr t = map f (Fr t) *)
    + assert (Fr t = map f (Fr t)) as A. 2: apply A.

      (* Again by transitivity ... *)
      apply eq_trans with (map id (Fr t)).

      (* ... it is sufficient to show firstly that Fr t = map id (Fr t) *)
      * assert (Fr t = map id (Fr t)) as A. 2: apply A.

        symmetry. apply map_id.

      (* ... and secondly that map id (Fr t) = map f (Fr t) ... *)
      * assert (map id (Fr t) = map f (Fr t)) as A. 2: apply A.

        (* ... which is the case ... *)
        apply coincide_map.

        (* ... provided we show that id and f coincide on Fr t  *)
        assert (coincide (Fr t) id f) as A. 2: apply A.

        (* So let u be a free variable of t *)
        intros u H2.

        (* We need to show that id u = f u *)
        assert (id u = f u) as A. 2: apply A.

        destruct H1 as [H1 H3]. symmetry. apply H3, H2.

    + assert (map f (Fr t) = Fr (fmap f t)) as A. 2: apply A.

      symmetry. destruct H1 as [H1 H3]. 

      apply (valid_free v v e e f t).
        { apply H1. }
        { apply Sub_refl. }
Qed.

(* The binding variable does not matter when not free *) 
Lemma Alpha_not_free_bind : forall (v:Type) (e:Eq v) (t1:T v) (x y:v),
  ~ x :: Fr t1 -> ~ y :: Fr t1 -> Lam x t1 ~ Lam y t1. 
Proof.
  (* Let v be a Type with decidable equality e *)
  intros v e.

  (* Let t1 be a term and x y be variables *)
  intros t1 x y.

  (* We assume that x and y are not free variables of t1 *)
  intros Hx Hy.

  (* We need to distinguish two cases *)
  destruct (eqDec x y) as [H1|H1].

  (* First we assume that x = y *)
  - rewrite <- H1.

    (* We need to show that Lam x t1 ~ All x t1 *)
    assert (Lam x t1 ~ Lam x t1) as A. 2: apply A.

    (* which is true by reflexivity *)
    apply Cong_reflexive.
  
  (* Next we assume that x <> y *)
  -
    (* We need to show that Lam x t1 is alpha-equivalent to Lam y t1 *)
    assert (Lam x t1 ~ Lam y t1) as A. 2: apply A.

    (* By transitivity, it is sufficient to prove two equivalences *)
    apply Cong_transitive with (Lam y (fmap (y <:> x) t1)).

    (* First we need to show that Lam x t1 ~ Lam y (fmap (y <:> x) t1) *)
    + assert (Lam x t1 ~ Lam y (fmap (y <:> x) t1)) as A. 2: apply A.

      (* This is true by definition of alpha-equivalence *)
      constructor. constructor.

      (* since  we have x <> y *)
      * assert (x <> y) as A. 2: apply A. apply H1.

      (* and y is not free in t1 *)
      * assert (~ y :: Fr t1) as A. 2: apply A. apply Hy.

    (* Second we need to show that Lam y (fmap (y <:> x) t1) ~ Lam y t1 *)
    + assert (Lam y (fmap (y <:> x) t1) ~ Lam y t1) as A. 2: apply A.

      apply CongLam. apply Cong_symmetric.

      (* So it is sufficient to show that fmap (y <:> x) t1 ~ t1 *)
      assert (t1 ~ fmap (y <:> x) t1) as A. 2: apply A.
  
      (* Using lemma Alpha_admissible, it is sufficient to show *)
      apply Alpha_admissible.

      (* that (y <:> x) is admissible for t1 *) 
      assert (admissible (y <:> x) t1) as A. 2: apply A.

      (* which follows from lemma admissible_permute *)
      apply admissible_permute.

        (* and the hypothesis of x y not free in t1 *)
        * assert (~ x :: Fr t1) as A. 2: apply A. apply Hx. 
        * assert (~ y :: Fr t1) as A. 2: apply A. apply Hy.
Qed.

(* Alpha-equivalence is preserved by injective maps *)
Lemma Alpha_injective :
  forall (v w:Type) (e:Eq v) (e':Eq w) (f:v -> w) (t s:T v),
    injective f -> t ~ s -> fmap f t ~ fmap f s.
Proof.
  (* Let v w be types with respective decidable equality e e' *)
  intros v w e e'.

  (* Let f be a map from v to w and t s be terms *)
  intros f t s.

  (* We assume that f is injective *)
  intros HInj. assert (injective f) as A. apply HInj. clear A.

  (* We need to show the implication t ~ s -> fmap f t ~ fmap f s *)
  assert (t ~ s -> fmap f t ~ fmap f s) as A. 2: apply A.

  (* Define the relation r as r t s = fmap f t ~ fmap f s *)
  remember (fun (t s:T v) => fmap f t ~ fmap f s) as r eqn:Er.

  (* Then r t s = fmap f t ~ fmap f s *)
  assert (r t s = fmap f t ~ fmap f s) as E. rewrite Er. reflexivity.

  (* So we need to show the implication t ~ s -> r t s for all t s *)
  rewrite <- E. clear E. revert s. revert t.
  assert (forall (t s:T v), t ~ s -> r t s) as A. 2: apply A.

  (* In other words, we need to show thw inclusion ~ <= r *)
  rewrite <- incl_charac.
  assert (Alpha <= r) as A. 2: apply A.

  (* Alpha being the smallest congruence on T v which contains Alpha0 *)
  apply Cong_smallest.

  (* It is sufficient first show that r is a congruence on T v *)
  - assert (congruence r) as A. 2: apply A. 

    (* which follows from Lemma fmap_congruence *)
    rewrite Er. apply fmap_congruence.

    (* together with the fact that alpha-equivalence is itself a congruence *)
    assert (congruence Alpha) as A. 2: apply A.

    (* which is true since Alpha is the congruence generated by Alpha0 *)
    apply Cong_congruence.

  (* and second to show that r contains Alpha0 *)
  - assert (Alpha0 <= r) as A. 2: apply A.

    (* So let x y be variables and t1 be a term *)
    rewrite incl_charac.
    intros t' s' H. destruct H as [x y t1 H3 H4]. 

    (* such that x <> y *)
    assert (x <> y) as A. apply H3. clear A. 

    (* and y is not free in t1 *)
    assert (~ y :: Fr t1) as A. apply H4. clear A.

    (* Define t = Lam x t1 *)
    remember (Lam x t1) as t eqn:Et.

    (* Define q = Lam y (fmap (y <:> x) t1) *)
    remember (Lam y (fmap (y <:> x) t1)) as s eqn:Es.

    (* Then we simply need to show that r t s holds *)
    assert (r t s) as A. 2: apply A.

    (* or in other words that fmap f t ~ fmap f s *)
    rewrite Er.
    assert (fmap f t ~ fmap f s) as A. 2: apply A.

    (* It is sufficient to show that Alpha0 (fmap f t) (fmap f s) *)
    apply CongBase.
    assert (Alpha0 (fmap f t) (fmap f s)) as A. 2: apply A.

    (* So it is sufficient to show the existence of t1' : T w
       and x' y' : w with x' <> y' and y' not free in t1' such that
       fmap f t = Lam x' t1' and fmap f s = Lam y' (fmap (y'<:>x') t1') *)
    
    (* Define t1' = fmap f t1 *)
    remember (fmap f t1) as t1' eqn:Et1'.
    
    (* Define x' = f x *)
    remember (f x) as x' eqn:Ex'.

    (* Define y' = f y *)
    remember (f y) as y' eqn:Ey'.

    (* Then we do have fmap f t = Lam x' t1' *)
    assert (fmap f t = Lam x' t1') as E1.
      { rewrite Et, Ex', Et1'. reflexivity. }

    (* and fmap f s = Lam y' (fmap <y':x'> t1') *)
    assert (fmap f s = Lam y' (fmap (y'<:>x') t1')) as E2.
      { rewrite Es, Ex', Ey', Et1'. simpl.
        rewrite <- fmap_comp', <- fmap_comp'.
        rewrite <- (permute_comp v w e e'). 
        reflexivity. 
        apply HInj. (* f is injective *)
      }

    (* we also have x' <> y' *)
    assert (x' <> y') as HNeq.
      { rewrite Ex', Ey'. intro H. apply HInj in H. contradiction. } 

    (* and y' is not free in t1' *)
    assert (~ y' :: Fr t1') as HFree.
    { rewrite Et1'. rewrite (free_inj v w e e'). 
      2: apply injective_injective_on, HInj.
      intro HFree. apply in_map_iff in HFree. 
      destruct HFree as [u [H1 H2]].
      rewrite Ey' in H1. apply HInj in H1. subst. 
      contradiction.
    }

    (* which allows us to conclude *)
    rewrite E1,E2. constructor.
      { apply HNeq. }
      { apply HFree. }
Qed.

(* Almost alpha-equivalence. Will be shown to be the same *)
Inductive AlmostAlpha (v:Type) (e:Eq v) : T v -> T v -> Prop :=
| AVar : forall (x:v), AlmostAlpha v e (Var x) (Var x)  
| AApp : forall (t1 t2 s1 s2:T v),
    t1 ~ s1 ->
    t2 ~ s2 ->
    AlmostAlpha v e (App t1 t2) (App s1 s2)
|ALamx : forall (x:v) (t1 s1:T v),
  t1 ~ s1 ->
  AlmostAlpha v e (Lam x t1) (Lam x s1)
| ALamxy : forall (x y:v) (t1 s1:T v),
  x <> y                  ->
  s1 ~ fmap (y <:> x) t1  ->
  ~ y :: Fr t1            ->
  AlmostAlpha v e (Lam x t1) (Lam y s1)
.

Arguments AlmostAlpha {v} {e}.

Notation "t :~: s" := (AlmostAlpha t s)
    (at level 60, no associativity) : Lam_Alpha_scope.

Open Scope Lam_Alpha_scope.

Lemma almostAppRev : forall (v:Type) (e:Eq v) (t1 t2 s:T v),
  App t1 t2 :~: s -> exists (s1 s2: T v),
    (t1 ~ s1) /\ (t2 ~ s2) /\ (s = App s1 s2).
Proof.
  (* Let v be a type with decidable equality e *)
  intros v e.

  (* Let t1 t2 s be formulas *)
  intros t1 t2 s.

  (* Define t = App t1 t2 *)
  remember (App t1 t2) as t eqn:Et.

  (* We assume that t is almost alpha-equivalent to s *)
  intro Haeq. assert (t :~: s) as A. apply Haeq. clear A.

  (* So we want to show that for all t1 t2 such that t = App t1 t2 ... *)
  revert t1 t2 Et.

  (* Case analysis on the assumption Haeq *)
  destruct Haeq as [x|t1' t2' s1 s2 H1 H2|x t1' s1|x y t1' s1 H1 H2 H3];
  intros t1 t2 Et.  
  
  (* Case t = s = Var x: Var x = App t1 t2 is a contradiction *)
  - inversion Et.

  (* Case t = App p1' p2' , s = App s1 s2 *)
  - inversion Et. subst. exists s1, s2. split.
      { assert (t1 ~ s1) as A. 2: apply A. apply H1. }
      { split.
        { assert (t2 ~ s2) as A. 2: apply A. apply H2. }
        { assert (App s1 s2 = App s1 s2) as A. 2: apply A. reflexivity. }
      } 
  (* Case t = Lam x t1' and s = Lam x s1: another contradiction *) 
  - inversion Et.
      
  (* Case t = Lam x t1' and s = Lam y s1: another contradiction *) 
  - inversion Et.
Qed.
