Require Import List.

Require Import Logic.Class.Eq.

Require Import Logic.Rel.R.
Require Import Logic.Rel.Include.

Require Import Logic.Func.Permute.
Require Import Logic.Func.Identity.
Require Import Logic.Func.Injective.
Require Import Logic.Func.Composition.

Require Import Logic.List.In.
Require Import Logic.List.Remove.
Require Import Logic.List.Append.
Require Import Logic.List.InjectiveOn.

Require Import Logic.Lam.Free.
Require Import Logic.Lam.Valid.
Require Import Logic.Lam.Syntax.
Require Import Logic.Lam.Functor.
Require Import Logic.Lam.Variable.
Require Import Logic.Lam.Congruence.
Require Import Logic.Lam.Admissible.

(* Generator of alpha-equivalence.                                              *)
(* We wish to formally define alpha-equivalence as the smallest congruence      *)
(* contaning all ordered pairs below. Note that we are using the permutation    *)
(* y <:> x rather than the substitution (y // x) and we allow the variable y    *)
(* to be a variable of t1 as long as it is not free. This seemingly unusual     *)
(* choice is to make sure we obtain a definition of alpha-equivalence which     *)
(* works equally well for a finite or infinite variable type v. Otherwise, we   *)
(* would obtain a congruence which is strictly stronger than alpha-equivalence  *)
(* when v is finite. See the StrongAlpha module for details.                    *)
Inductive Alpha0 (v:Type) (e:Eq v) : T v -> T v -> Prop :=
| mkAlpha0: forall (x y:v) (t1:T v), 
    x <> y       -> 
    ~ y :: Fr t1 ->
    Alpha0 v e (Lam x t1) (Lam y (fmap (y <:> x) t1)) 
.

Arguments Alpha0 {v} {e}.
Arguments mkAlpha0 {v} {e}.

(* The alpha-equivalence relation is the congruence generated by Alph0.         *)
Definition Alpha (v:Type) (e:Eq v) : T v -> T v -> Prop := 
    Cong (@Alpha0 v e).

Arguments Alpha {v} {e}.

Notation "t ~ s" := (Alpha t s)
    (at level 60, no associativity) : Lam_Alpha_scope.

Open Scope Lam_Alpha_scope.

(* Admissible substitutions do not change alpha-equivalence classes.            *)
Lemma Alpha_admissible : forall (v:Type) (e:Eq v) (t:T v) (f:v -> v),
  admissible f t -> t ~ fmap f t.
Proof.
  intros v e.
  induction t as [x|t1 IH1 t2 IH2|x t1 IH1]; 
  intros f [H1 H2]; simpl; simpl in H2.

  (* case t = Var x *)
  - assert (f x = x) as E1. { apply H2. left. reflexivity. }
    rewrite E1. apply Cong_reflexive.

  (* case t = App t1 t2 *)
  - rewrite valid_app in H1; destruct H1 as [H1 H3].

    assert (t1 ~ fmap f t1) as E1.
      { apply IH1. unfold admissible. split.
        { assumption. }
        { intros x H4. apply H2, app_charac. left. assumption. }}

    assert (t2 ~ fmap f t2) as E2.
      { apply IH2. unfold admissible. split.
        { assumption. }
        { intros x H4. apply H2, app_charac. right. assumption. }}

    apply CongApp; assumption. 

  (* case t = Lam x t1 *)
  - rewrite valid_lam in H1. destruct H1 as [H3 H4].
    destruct (eqDec (f x) x) as [H5|H5].

    + (* f x = x *)
      assert (t1 ~ fmap f t1) as E1.
        { apply IH1. unfold admissible. split.
          { assumption. }
          { intros y H6.
            assert (f y = y) as E1.
              { destruct (eqDec x y) as [H7|H7].
                { (* x = y  *)
                  rewrite <- H7. assumption. }
                { (* x <> y *)
                  apply H2, remove_charac. split; assumption. }}
           assumption. }} 
      rewrite H5. apply CongLam. assumption.
      
    + (* f x <> x *)
      remember (f x) as y eqn:H6.

      assert (Lam x t1 ~ Lam y (fmap f t1)) as E.
        { remember ((y <:> x) ; f) as g eqn:H7.
          remember (fmap g t1) as s1 eqn:H8. 

          assert (f = (y <:> x) ; g) as E1.
            { rewrite H7. rewrite comp_assoc, permute_involution.
              symmetry. apply comp_id_left. }

          assert (fmap f t1 = fmap (y <:> x) s1) as E2.
            { rewrite H8, <- fmap_comp', <- E1. reflexivity. }

          rewrite E2.

          assert (Lam x t1 ~ Lam y (fmap (y <:> x) s1)) as E3.
            { assert (admissible g t1) as E8. 
                { unfold admissible. split.
                   { rewrite H7. rewrite <- valid_compose. split.
                    { apply H3. (* why is the assumption tactic failing here *) }
                    { apply valid_inj, injective_injective_on. 
                      apply permute_injective. }}
                { intros u H10. destruct (eqDec u x) as [H11|H11].
                    { subst. unfold comp. apply permute_app_left. }
                    { rewrite H7. unfold comp. 
                      assert (f u = u) as H12.
                        { apply H2. apply remove_charac. split.
                            { assumption. }
                            { apply not_eq_sym.  assumption. }}
                      rewrite H12. apply permute_app_diff. 
                        { intros H13. apply H4 with u. 
                          { simpl. apply remove_charac. split.
                            { assumption. }
                            { apply not_eq_sym. assumption. }}
                          { rewrite H12. symmetry. assumption. }}
                        { assumption. }}}}

              assert (~ y :: Fr s1) as E4.
                { rewrite H8. intros H9. apply (free_fmap v v e) in H9.
                  apply in_map_iff in H9. destruct H9 as [u [H9 H10]].
                  unfold admissible in E8. destruct E8 as [H11 H12]. 
        
                  assert (g u = u) as H13. { apply H12. assumption. }

                  assert (y :: Fr t1) as H14. { rewrite <- H9, H13. assumption. }
              
                  assert (y :: Fr (Lam x t1)) as H15.
                    { simpl. apply remove_charac. split.
                      { assumption. }
                      { apply not_eq_sym. assumption. }} 

                  assert (f y = y) as H17. { apply H2. assumption. }

                  assert (f x <> f y) as H18. 
                    { rewrite <- H6. apply H4. assumption. }

                  assert (f x <> y) as H19. { rewrite <- H17. assumption. }
  
                  apply H19. symmetry. assumption. }

              assert (Lam x s1 ~ Lam y (fmap (y <:> x) s1)) as E5.
                { constructor. constructor.
                  { intros H9. apply H5. symmetry. assumption. }
                  { assumption. }}

              assert (Lam x t1 ~ Lam x s1) as E6.
                { assert (t1 ~ s1) as E7. { rewrite H8. apply IH1. apply E8. }
                  apply Cong_congruent, E7. }

              apply Cong_transitive with (Lam x s1); assumption. }
          apply E3. }
      apply E.
Qed.

(* This is a relation which is larger than Alpha0 but a lot simpler. As we      *)
(* shall see, it is also a generator of the alpha-equivalence congruence.       *)
Inductive Alpha1 (v:Type) (e:Eq v) : T v -> T v -> Prop :=
| mkAlpha1: forall (t:T v) (f:v -> v), admissible f t -> Alpha1 v e t (fmap f t)
.

Arguments Alpha1 {v} {e}.
Arguments mkAlpha1 {v} {e}.

(* Alpha-equivalence is also the congruence generated by Alpha1.                *)
Lemma Alpha_admissible_gen : forall (v:Type) (e:Eq v), Alpha = Cong Alpha1.
Proof.
  intros v e.  
  remember (Cong Alpha1) as r eqn:E1.

  assert (Alpha <= r) as A1.
    { assert (Alpha0 <= r) as A2.
        { apply incl_charac. intros t s H1. destruct H1 as [x y t1 H1 H2].
          remember (Lam x t1) as t eqn:E2.
          remember (Lam y (fmap (y <:> x) t1)) as s eqn:E3.

          assert (Alpha1 t s) as A3.
            { remember (y <:> x) as f eqn:E4.

              assert (s = fmap f t) as A4.
                { rewrite E2, E3. simpl.

                  assert (f x = y) as A5. { rewrite E4. apply permute_app_right. }
                  rewrite A5. reflexivity. }

              rewrite A4. constructor.  

              assert (admissible f t) as A6.
                { unfold admissible. split. 

                    { assert (valid f t) as A7.
                        { apply valid_inj, injective_injective_on.

                          assert (injective f) as A8.
                            { rewrite E4. apply permute_injective. }
                          apply A8. }

                      apply A7. }

                    { assert (forall (u:v), u :: Fr t -> f u = u) as A9.
                        { intros u H3.

                          assert (u <> x) as A10.
                            { rewrite E2 in H3. simpl in H3. 
                              apply remove_charac in H3.
                              destruct H3 as [H3 H4]. apply not_eq_sym.
                              assumption. }
  
                          assert (u <> y) as A11.
                            { assert (u :: Fr t1) as A12.
                                { rewrite E2 in H3. simpl in H3.
                                  apply remove_charac in H3.
                                  destruct H3 as [H3 H4]. assumption. }

                              intros H4. rewrite H4 in A12. contradiction. } 
 
                          rewrite E4. apply permute_app_diff; assumption. }


                      apply A9. } }

              apply A6. }

          rewrite E1. constructor. apply A3. } 

      unfold Alpha. apply Cong_smallest.
        { assert (congruence r) as A13.
            { rewrite E1. apply Cong_congruence. }

          apply A13. }

        { apply A2. } }

  assert (r <= Alpha) as A14.
    { assert (Alpha1 <= Alpha) as A15.
        { apply incl_charac. intros t s H5. destruct H5 as [t f H5].
          apply Alpha_admissible. assumption. }

      rewrite E1. apply Cong_smallest.
        { assert (congruence Alpha) as A16.
            { unfold Alpha. apply Cong_congruence. }

          apply A16. }

        { apply A15. } }

  apply incl_anti.
    { apply A1. }
    { apply A14. }
Qed.
