Require Import List.

Require Import Logic.Class.Eq.

Require Import Logic.Rel.R.
Require Import Logic.Rel.Include.

Require Import Logic.Func.Permute.
Require Import Logic.Func.Identity.
Require Import Logic.Func.Injective.
Require Import Logic.Func.Composition.

Require Import Logic.List.In.
Require Import Logic.List.Remove.
Require Import Logic.List.Append.
Require Import Logic.List.InjectiveOn.

Require Import Logic.Fol.Free.
Require Import Logic.Fol.Valid.
Require Import Logic.Fol.Syntax.
Require Import Logic.Fol.Functor.
Require Import Logic.Fol.Variable.
Require Import Logic.Fol.Congruence.
Require Import Logic.Fol.Admissible.

(* Generator of alpha-equivalence.                                              *)
(* We wish to formally define alpha-equivalence as the smallest congruence      *)
(* contaning all ordered pairs below. Note that we are using the permutation    *)
(* y <:> x rather than the substitution (y // x) and we allow the variable y    *)
(* to be a variable of p1 as long as it is not free. This seemingly unusual     *)
(* choice is to make sure we obtain a definition of alpha-equivalence which     *)
(* works equally well for a finite or infinite variable type v. Otherwise, we   *)
(* would obtain a congruence which is strictly stronger than alpha-equivalence  *)
(* when v is finite. See the StrongAlpha module for details.                    *)
Inductive Alpha0 (v:Type) (e:Eq v) : P v -> P v -> Prop :=
| mkAlpha0: forall (x y:v) (p1:P v), 
    x <> y       -> 
    ~ y :: Fr p1 ->
    Alpha0 v e (All x p1) (All y (fmap (y <:> x) p1)) 
.

Arguments Alpha0 {v} {e}.
Arguments mkAlpha0 {v} {e}.

(* The alpha-equivalence relation is the congruence generated by Alph0.         *)
Definition Alpha (v:Type) (e:Eq v) : P v -> P v -> Prop := 
    Cong (@Alpha0 v e).

Arguments Alpha {v} {e}.

Notation "p ~ q" := (Alpha p q)
    (at level 60, no associativity) : Fol_Alpha_scope.

Open Scope Fol_Alpha_scope.

(* Admissible substitutions do not change alpha-equivalence classes.            *)
Lemma Alpha_admissible : forall (v:Type) (e:Eq v) (p:P v) (f:v -> v),
  admissible f p -> p ~ fmap f p.
Proof.
  intros v e.
  induction p as [|x y|p1 IH1 p2 IH2|x p1 IH1]; 
  intros f [H1 H2]; simpl; simpl in H2.

  (* case p = Bot *)
  - apply Cong_reflexive.

  (* case p = Elem x y *)
  - assert (f x = x) as E1. { apply H2. left. reflexivity. }
    assert (f y = y) as E2. { apply H2. right. left. reflexivity. }
    rewrite E1, E2. apply Cong_reflexive.

  (* case p = Imp p1 p2 *)
  - rewrite valid_imp in H1; destruct H1 as [H1 H3].

    assert (p1 ~ fmap f p1) as E1.
      { apply IH1. unfold admissible. split.
        { assumption. }
        { intros x H4. apply H2, app_charac. left. assumption. }}

    assert (p2 ~ fmap f p2) as E2.
      { apply IH2. unfold admissible. split.
        { assumption. }
        { intros x H4. apply H2, app_charac. right. assumption. }}

    apply CongImp; assumption. 

  (* case p = All x p1 *)
  - rewrite valid_all in H1. destruct H1 as [H3 H4].
    destruct (eqDec (f x) x) as [H5|H5].

    + (* f x = x *)
      assert (p1 ~ fmap f p1) as E1.
        { apply IH1. unfold admissible. split.
          { assumption. }
          { intros y H6.
            assert (f y = y) as E1.
              { destruct (eqDec x y) as [H7|H7].
                { (* x = y  *)
                  rewrite <- H7. assumption. }
                { (* x <> y *)
                  apply H2, remove_charac. split; assumption. }}
           assumption. }} 
      rewrite H5. apply CongAll. assumption.

    + (* f x <> x *)
      remember (f x) as y eqn:H6.

      assert (All x p1 ~ All y (fmap f p1)) as E.
        { remember ((y <:> x) ; f) as g eqn:H7.
          remember (fmap g p1) as q1 eqn:H8. 

          assert (f = (y <:> x) ; g) as E1.
            { rewrite H7. rewrite comp_assoc, permute_involution.
              symmetry. apply comp_id_left. }

          assert (fmap f p1 = fmap (y <:> x) q1) as E2.
            { rewrite H8, <- fmap_comp', <- E1. reflexivity. }

          rewrite E2.

          assert (All x p1 ~ All y (fmap (y <:> x) q1)) as E3.
            { assert (admissible g p1) as E8. 
                { unfold admissible. split.
                  { rewrite H7. rewrite <- valid_compose. split.
                    { apply H3. (* why is the assumption tactic failing here *) }
                    { apply valid_inj, injective_injective_on. 
                      apply permute_injective. }}
                  { intros u H10. destruct (eqDec u x) as [H11|H11].
                    { subst. unfold comp. apply permute_app_left. }
                    { rewrite H7. unfold comp. 
                      assert (f u = u) as H12.
                        { apply H2. apply remove_charac. split.
                            { assumption. }
                            { apply not_eq_sym.  assumption. }}
                      rewrite H12. apply permute_app_diff. 
                        { intros H13. apply H4 with u. 
                          { simpl. apply remove_charac. split.
                            { assumption. }
                            { apply not_eq_sym. assumption. }}
                          { rewrite H12. symmetry. assumption. }}
                        { assumption. }}}}

              assert (~ y :: Fr q1) as E4.
                { rewrite H8. intros H9. apply (free_fmap v v e) in H9.
                  apply in_map_iff in H9. destruct H9 as [u [H9 H10]].
                  unfold admissible in E8. destruct E8 as [H11 H12]. 

                  assert (g u = u) as H13. { apply H12. assumption. }

                  assert (y :: Fr p1) as H14. { rewrite <- H9, H13. assumption. }

                  assert (y :: Fr (All x p1)) as H15.
                    { simpl. apply remove_charac. split.
                      { assumption. }
                      { apply not_eq_sym. assumption. }} 

                  assert (f y = y) as H17. { apply H2. assumption. }

                  assert (f x <> f y) as H18. 
                    { rewrite <- H6. apply H4. assumption. }

                  assert (f x <> y) as H19. { rewrite <- H17. assumption. }

                  apply H19. symmetry. assumption. }

              assert (All x q1 ~ All y (fmap (y <:> x) q1)) as E5.
                { constructor. constructor.
                  { apply not_eq_sym. assumption. }
                  { assumption. }}

              assert (All x p1 ~ All x q1) as E6.
                { assert (p1 ~ q1) as E7. { rewrite H8. apply IH1. apply E8. }
                  apply Cong_congruent, E7. }

              apply Cong_transitive with (All x q1); assumption. }
          apply E3. }
      apply E.
Qed.

(* This is a relation which is larger than Alpha0 but a lot simpler. As we      *)
(* shall see, it is also a generator of the alpha-equivalence congruence.       *)
Inductive Alpha1 (v:Type) (e:Eq v) : P v -> P v -> Prop :=
| mkAlpha1: forall (p:P v) (f:v -> v), admissible f p -> Alpha1 v e p (fmap f p)
.

Arguments Alpha1 {v} {e}.
Arguments mkAlpha1 {v} {e}.

(* Alpha-equivalence is also the congruence generated by Alpha1.                *)
Lemma Alpha_admissible_gen : forall (v:Type) (e:Eq v), Alpha = Cong Alpha1.
Proof.
  (* Let v be a Type with decidable equality e  *)
  intros v e.
  
  (* Define r  *)
  remember (Cong Alpha1) as r eqn:E1.

  (* We need to show that Alpha = r *)
  assert (Alpha = r) as A. 2: apply A.

  (* We do so with a double inclusion argument *)
  apply incl_anti.

  (* First we show that Alpha <= r  *)
  - assert (Alpha <= r) as A. 2: apply A.

    (* We argue that Alpha is the smallest congruence containing Alpha0 *)
    unfold Alpha. apply Cong_smallest.

      (* So we need to show that r is a congruence  *)
      + assert (congruence r) as A. 2: apply A.
        
        rewrite E1. apply Cong_congruence.

      (* And we need to show that r contains Alpha0 *)
      + assert (Alpha0 <= r) as A. 2: apply A.

        (* So let x y and p1 such that x <> y and ~ y :: Fr p1  *)
        apply incl_charac. intros p q H1. destruct H1 as [x y p1 H1 H2].

        (* Define p *)
        remember (All x p1) as p eqn:E2.

        (* Define q *)
        remember (All y (fmap (y <:> x) p1)) as q eqn:E3.

        (* Define f *)
        remember (y <:> x) as f eqn:E4.

        (* We need to show that (p,q) :: r  *)
        assert (r p q) as A. 2: apply A.

        (* i.e. that (p.q) belongs to the congruence generated by Alpha1  *)
        rewrite E1. 
        
        (* We argue that (p,q) actually belongs to the generator itself *)
        constructor.

        (* So we need to show that (p,q) belongs to Alpha1  *)
        assert (Alpha1 p q) as A. 2: apply A.

        (* However, q is in fact q = fmap f p *)
        assert (q = fmap f p) as A.
          { rewrite E2, E3. simpl.
            assert (f x = y) as A5. 2: rewrite A5; reflexivity.
            rewrite E4. apply permute_app_right.
          }

        (* So we need to show that (p, fmap f p) lies in Alpha1 *)
        rewrite A. clear A. 
          
        (* which is true by definition... *)
        constructor.  
    
        (* ... provided we show that f is admissible for p  *)
        assert (admissible f p) as A. 2: apply A.
        
        (* Given the definition of an admissible substitution *)
        unfold admissible. split. 

          (* First we need to show that f is valid for p *)
          * assert (valid f p) as A. 2: apply A.
            
            (* It is sufficient to show that f is injective on (var p) *)
            apply valid_inj.
            
            (* It is sufficient to show that f is injective *)
            apply injective_injective_on.

            (* So we now prove that f is injective *)
            assert (injective f) as A. 2: apply A. 
            
            (* However, f is the permutation mapping (y <:> x)  *) 
            rewrite E4. 
            
            (* it is therefore injective  *)
            apply permute_injective.
         

          (* And furthermore that free variables are invariant by f *)
          * assert (forall (u:v), u :: Fr p -> f u = u) as A. 2: apply A.
            
            (* So let u with u :: Fr p  *) 
            intros u H3.
            
            (* We need to show that f u = u *)
            assert (f u = u) as A. 2: apply A.

            (* Given that f is the permutation mapping (y <:> x) ...  *)
            rewrite E4.

            (* ... it is sufficient to show that u <> x and u <> y *)
            apply permute_app_diff. 

              (* First we show that u <> y  *)
              { assert (u <> y) as A. 2: apply A.

                (* Since u :: Fr p, we have u :: Fr p1  *)
                assert (u :: Fr p1) as A.
                  { rewrite E2 in H3. simpl in H3.
                    apply remove_charac in H3.
                    destruct H3 as [H3 H4]. assumption. 
                  }
                
                (* So if we assume that u = y ... *)
                intros H4. 

                (* ... we obtain y :: Fr p1 which is a contradiction  *)
                rewrite H4 in A. contradiction. 
              }

              (* We now show that u <> x  *)
              { assert (u <> x) as A. 2: apply A.

                (* This is the case since u is free in p = All x p1 *)
                rewrite E2 in H3. simpl in H3. 
                apply remove_charac in H3.
                destruct H3 as [H3 H4]. apply not_eq_sym.
                assumption.

              } 
          
  (* We now show that r <= Alpha  *)
  - assert (r <= Alpha) as A. 2: apply A.
    
    (* We argue that r is the smallest congruence containing Alpha1 *)
    rewrite E1. apply Cong_smallest.

    (* So we need to show that Alpha is a congruence  *)
    + assert (congruence Alpha) as A. 2: apply A.
      
      (* Given that Alpha is the congruence generated by Alpha0 ... *)
      unfold Alpha. 
        
      (* ... it is indeed a congruence  *)
      apply Cong_congruence.
 
    (* And we need to show that Alpha contains Alpha1 *)
    + assert (Alpha1 <= Alpha) as A. 2: apply A.
      
      (* So let p and f : v -> v such that f is admissible *) 
      apply incl_charac. intros p q H5. destruct H5 as [p f H5].

      (* We need to show that p is alpha-equivalent to fmap f p  *)
      assert (p ~ fmap f p) as A. 2: apply A. 

      (* This is the case, provided f is admissible ... *)
      apply Alpha_admissible. 
      
      (* ... which is true by assumption *)
      assumption. 
   
Qed.

(*
(* Not following pdf to obtain stronger result of equality as lists.            *)
(* Two alpha-equivalent formulas have the same free variables.                  *)
Lemma Alpha_free : forall (v:Type) (e:Eq v) (p q:P v), 
    p ~ q -> Fr p = Fr q.
Proof.
  intros v e.  
  remember (fun (p q:P v) => Fr p = Fr q) as r eqn:E1.
  apply incl_charac. rewrite <- E1. 

  (* We simply need to show that Alpha <= r *)
  assert (Alpha <= r) as A1. 2 : apply A1. 


Show.
*)
