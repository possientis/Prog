Require Import List.

Require Import Logic.Class.Eq.

Require Import Logic.Rel.R.
Require Import Logic.Rel.Include.

Require Import Logic.Func.Permute.
Require Import Logic.Func.Identity.
Require Import Logic.Func.Injective.
Require Import Logic.Func.Composition.

Require Import Logic.List.In.
Require Import Logic.List.Remove.
Require Import Logic.List.Append.
Require Import Logic.List.Coincide.
Require Import Logic.List.InjectiveOn.

Require Import Logic.Fol.Free.
Require Import Logic.Fol.Valid.
Require Import Logic.Fol.Syntax.
Require Import Logic.Fol.Functor.
Require Import Logic.Fol.Variable.
Require Import Logic.Fol.Congruence.
Require Import Logic.Fol.Subformula.
Require Import Logic.Fol.Admissible.

Declare Scope Fol_Alpha_scope.

(* Generator of alpha-equivalence.                                              *)
(* We wish to formally define alpha-equivalence as the smallest congruence      *)
(* contaning all ordered pairs below. Note that we are using the permutation    *)
(* y <:> x rather than the substitution (y // x) and we allow the variable y    *)
(* to be a variable of p1 as long as it is not free. This seemingly unusual     *)
(* choice is to make sure we obtain a definition of alpha-equivalence which     *)
(* works equally well for a finite or infinite variable type v. Otherwise, we   *)
(* would obtain a congruence which is strictly stronger than alpha-equivalence  *)
(* when v is finite. See the StrongAlpha module for details.                    *)
Inductive Alpha0 (v:Type) (e:Eq v) : P v -> P v -> Prop :=
| mkAlpha0: forall (x y:v) (p1:P v), 
    x <> y       -> 
    ~ y :: Fr p1 ->
    Alpha0 v e (All x p1) (All y (fmap (y <:> x) p1)) 
.

Arguments Alpha0 {v} {e}.
Arguments mkAlpha0 {v} {e}.

(* The alpha-equivalence relation is the congruence generated by Alph0.         *)
Definition Alpha (v:Type) (e:Eq v) : P v -> P v -> Prop := 
    Cong (@Alpha0 v e).

Arguments Alpha {v} {e}.

Notation "p ~ q" := (Alpha p q)
    (at level 60, no associativity) : Fol_Alpha_scope.

Open Scope Fol_Alpha_scope.

(* Admissible substitutions do not change alpha-equivalence classes.            *)
Lemma Alpha_admissible : forall (v:Type) (e:Eq v) (p:P v) (f:v -> v),
  admissible f p -> p ~ fmap f p.
Proof.
  (* Let v be a Type with decidable equality e  *)
  intros v e.

  (* We prove the lemma with an induction argument on p *)
  induction p as [|x y|p1 IH1 p2 IH2|x p1 IH1]; 

  (* In each case we assume f:v -> v is admissible for p *)
  intros f H1.

  (* case p = Bot *)
  - assert (Bot ~ Bot) as A. 2: apply A.

    apply Cong_reflexive.

  (* case p = Elem x y *)
  - assert (Elem x y ~ Elem (f x) (f y)) as A. 2: apply A.

    assert (f x = x) as A1. 
    { apply admissible_free with (Elem x y).
      - apply H1.
      - left. reflexivity.
    }
    
    assert (f y = y) as A2. 
    { apply admissible_free with (Elem x y).
      - apply H1. 
      - right. left. reflexivity.
    }
      
    rewrite A1, A2. 

    apply Cong_reflexive.

  (* case p = Imp p1 p2 *)
  - assert (Imp p1 p2 ~ Imp (fmap f p1) (fmap f p2)) as A. 2: apply A. 

    (* Note that f being admissible for Imp p1 p2  ... *)
    apply admissible_imp in H1. destruct H1 as [H1 H2].
    
    (* ... it is admissible for p1 ... *)
    assert (admissible f p1) as A. apply H1. clear A.

    (* ... and it is admissible for p2 *)
    assert (admissible f p2) as A. apply H2. clear A.

    (* We argue that alpha-equivalence is a congruence  *)
    apply CongImp.

    (* So we need to prove that p1 ~ fmap f p1  *)
    + assert (p1 ~ fmap f p1) as A. 2: apply A. 
  
      (* This follows from the induction hypothesis ... *)
      apply IH1. 

      (* ... provided we show that f is admissible for p1 ... *)
      assert (admissible f p1) as A. 2: apply A.
    
      (* ... which we know is true  *) 
      apply H1.

    (* We need to prove similarly that p2 ~ fmap f p2  *)
    + assert (p2 ~ fmap f p2) as A. 2: apply A.

      (* This follows from the induction hypothesis ... *)
      apply IH2.

      (* ... provided we show that f is admissible for p2 ... *)
      assert (admissible f p2) as A. 2: apply A.

      (* ... which we know is true *)
      apply H2.

  (* case p = All x p1 *)
  - assert (All x p1 ~ All (f x) (fmap f p1)) as A. 2: apply A. 
   
    (* Note that f being admissible for All x p1 ... *)
    destruct H1 as [H1 H3]. apply valid_all in H1. destruct H1 as [H1 H2].

    (* ... it is valid for p1 ... *)
    assert (valid f p1) as A. apply H1. clear A.

    (* ... we have f x <> f y for any y free in All x p1  ... *)
    assert (forall (y:v), y :: Fr (All x p1)->f x <> f y) as A. apply H2. clear A.

    (* ... and we have f y = y for any y free in All x p1 *)
    assert (forall (y:v), y :: Fr (All x p1) -> f y = y) as A. apply H3. clear A.
 
    (* We carry out the proof by distinguishing two cases *)
    destruct (eqDec (f x) x) as [H4|H4].

    + (* First we assume that f x = x *)

      (* Given that f x = x *)
      rewrite H4.

      (* We need to show that All x p1 ~ All x (fmap f p1)  *)
      assert (All x p1 ~ All x (fmap f p1)) as A. 2: apply A.

      (* Alpha-equivalence being a congruence ... *)
      apply CongAll.

      (* ... we simply need to show that p1 ~ fmap f p1 *)
      assert (p1 ~ fmap f p1) as A. 2: apply A.

      (* This follows from the induction hypothesis ... *)
      apply IH1.

      (* ... provided we show that f is admissible for p1 *)
      assert (admissible f p1) as A. 2: apply A.

      (* Given the definition of an admissible mapping ... *)
      unfold admissible. split.

      (* ... we need to show that f is valid for p1 ... *)
      * assert (valid f p1) as A. 2: apply A.

        (* ... which is true as we have noted *)
        apply H1.

      (* ... and that free variables of p1 are invariant by f *)
      * assert (forall (u:v), u :: Fr p1 -> f u = u) as A. 2: apply A.

        (* So let u with u :: Fr p1 *)
        intros u H5. 
      
        (* We need to show that f u = u ... *) 
        assert (f u = u) as A. 2: apply A.

        (* We shall distinguish two cases *)
        destruct (eqDec x u) as [H6|H6].

        (* First we assume that x = u *)
        { rewrite <- H6.

          (* Then we need to show that f x = x ...  *)
          assert (f x = x) as A. 2: apply A.

          (* ... which we have assumed is true. *)
          apply H4.
        }

        (* Next we assume that x <> u *)
        { 
          (* Then f u = u follows from H3 ... *)
          apply H3.

          (* ... provided we show that u is free in All x p1  *) 
          assert (u :: Fr (All x p1)) as A. 2: apply A.
           
          simpl. apply remove_charac. split; assumption.
        }

    + (* Then we assume that f x <> x *)

      (* Define y *)
      remember (f x) as y eqn:E1.

      (* Define g *)
      remember ((y <:> x) ; f) as g eqn:E2.

      (* Define q1  *)
      remember (fmap g p1) as q1 eqn:E3. 

      (* So we need to show:  *)
      assert (All x p1 ~ All y (fmap f p1)) as A. 2: apply A.

      (* We claim that: *)
      assert (f = (y <:> x) ; g) as A1.
      { rewrite E2, comp_assoc, permute_involution. 
        symmetry. apply comp_id_left. 
      }
    
      (* And furthermore: *) 
      assert (fmap f p1 = fmap (y <:> x) q1) as A2.
      { rewrite E3, <- fmap_comp', <- A1. clear A1. reflexivity. 
      }

      (* We also claim that g is admissible for p1  *)
      assert (admissible g p1) as A3.
      { (* Given the definition of an admissible mapping ... *)
        unfold admissible. split.

        (* ... need need to show that g is valid for p1 *)
        - assert (valid g p1) as A. 2: apply A.
            
          (* Since g = (y <:> x) ; f  ... *)
          rewrite E2. 

          (* ... we need to show: *)
          assert (valid ((y <:> x) ; f) p1) as A. 2: apply A.

          (* and consequently ... *)
          rewrite <- valid_compose. split.

          (* ... we need to show that f is valid for p1 ... *)
          +  assert (valid f p1) as A. 2: apply A.
            
             (* ... we which know is true *)
             apply H1.

          (* ... and we need to show that (y <:> x) is valid for fmap f p1 ...*)
          + assert (valid (y <:> x) (fmap f p1)) as A. 2: apply A.

            (* ... which follows from the injectivity of pernutations *)
            apply valid_inj, injective_injective_on, permute_injective.

        (* ... and show that free variables of p1 are invariant by g  *)
        - assert (forall (u:v), u :: Fr p1 -> g u = u) as A. 2: apply A.

          (* so let u with u :: Fr p1 *)
          intros u H5. 

          (* We need to show that g u = u *)
          assert (g u = u) as A. 2: apply A.

          (* Given that g = (y <:> x) ... *)
          rewrite E2. unfold comp.

          (* ... amounts to showing that: *)
          assert ((y <:> x) (f u) = u) as A. 2: apply A.

          (* We shall distinguish two cases *)
          destruct (eqDec u x) as [H6|H6].

          * (* We first assume that u = x *)
           
            (* Given that u = x and y = f x ... *)
            rewrite H6, E1.

            (* ... we need to show that:  *)
            assert ((f x <:> x) (f x) = x) as A. 2: apply A.

            (* This is an immediate property of the permutation mapping *)
            apply permute_app_left.

          * (* We then assume that u <> x *)

            (* We claim that f u = u *)
            assert (f u = u) as A4.
            { (* This follows from H3 ... *)  
              apply H3. 

              (* ... provided we show that u is free in All x p1  *)
              assert (u :: Fr (All x p1)) as A. 2: apply A.

              simpl. apply remove_charac. split.

              (* So we need to show that u is free in p1 ...  *)
              - assert (u :: Fr p1) as A. 2: apply A.
                    
                apply H5.
              
              (* ... and that x <> u  *)
              - assert (x <> u) as A. 2: apply A.

                apply not_eq_sym, H6. 
            }             

            (* So given that f u = u ... *)
            rewrite A4.

            (* we need to show that:  *)
            assert ((y <:> x) u = u) as A. 2: apply A.

            (* Hence, it is sufficient to prove... *)
            apply permute_app_diff.

            (* ... that u <> y  *)
            { assert (u <> y) as A. 2: apply A.

              (* So suppose that u = y  *)
              intros H7.

              (* Then we obtain a contradiction by showing f u <> u *)
              assert (f u <> u) as A. 2: contradiction.

              (* Given that u = y ... *)
              apply not_eq_sym. rewrite H7 at 1.

              (* ... we need to show that y <> f u  *)
              assert (y <> f u) as A. 2: apply A. 

              (* This follows from H2 ... *)
              apply H2.

              (* ... provided we show that u is free in All x p1 *)
              assert (u :: Fr (All x p1)) as A. 2: apply A.
         
              simpl. apply remove_charac. split.

              (* So we need to show that u is free in p1 ...  *)
              - assert (u :: Fr p1) as A. 2: apply A.
                  
                apply H5.

              (* ... and that x <> u  *)
              - assert (x <> u) as A. 2: apply A. 
                
                apply not_eq_sym, H6. 
            }

            (* ... and u <> x  *)
            { assert (u <> x) as A. 2: apply A.
                  
              apply H6.
            }
      (* This completes the proof of the admissibility of g for p1  *)
      } 

      (* So we now need to show:  *)
      assert (All x p1 ~ All y (fmap f p1)) as A. 2: apply A.

      (* Given that fmap f p1 = fmap (y <:> x) q1 ... *)
      rewrite A2. clear A2.

      (* ... we need to show that:  *)
      assert (All x p1 ~ All y (fmap (y <:> x) q1)) as A. 2: apply A.

      (* Alpha-equivalence being a transitive relation ...  *)
      apply Cong_transitive with (All x q1).

      (* ... it is sufficient to show firstly that: *) 
      * assert (All x p1 ~ All x q1) as A. 2: apply A.

        (* Alpha-equivalence being a congruence ... *)
        apply Cong_congruent.

        (* ... it is sufficient to show that p1 ~ q1 *)
        assert (p1 ~ q1) as A. 2: apply A.

        (* Given that q1 = fmap g p1  *)
        rewrite E3.

        (* we need to show that p1 ~ fmap q p1 ... *)
        assert (p1 ~ fmap g p1) as A. 2: apply A.

        (* ... which follows from the induction hypothesis ... *)
        apply IH1.

        (* ... provided we show show that g is admissible for p1 ...  *)
        assert (admissible g p1) as A. 2: apply A.

        (* ... which we have already proven *)
        apply A3.

      (* ... and secondly that:  *)
      * assert (All x q1 ~ All y (fmap (y <:> x) q1)) as A. 2: apply A.

        (* We argue that the pair actually belongs to the generator Alpha0  *)
        constructor.

        (* So we need to show that: *)
        assert (Alpha0 (All x q1) (All y (fmap (y <:> x) q1))) as A. 2: apply A.

        (* This is true by definition ...  *)
        constructor.

        (* ... provided we show that x <> y ... *)
        { assert (x <> y) as A. 2: apply A. 
          
          (* ... which is true since with have assumed f x <> x *)
          apply not_eq_sym, H4.
        }

        (* ... and that y is not free in q1 *)
        { assert (~ y :: Fr q1) as A. 2: apply A. 

          (* Given that q1 = fmap g p1 ...  *)
          rewrite E3. 

          (* ... we need to show that y is not free in fmap g p1 *)
          assert (~ y :: Fr (fmap g p1)) as A. 2: apply A. 

          (* So suppose to the contrary that y is free in fmap g p1 *)
          intros H5. 

          (* We need to obtain a contradiction by showing y <> f x *)
          assert (y <> f x) as A. 2: contradiction.

          (* Since Fr (fmap g p1) <= map g (Fr p1), we have y :: map g (Fr p1)  *)
          apply (free_fmap v v e) in H5.

          (* So there exists u such that y = g u and u :: Fr p1 *)
          apply in_map_iff in H5. destruct H5 as [u [H5 H6]].

          (* Note that g is valid for p1 and g u = u for all u :: Fr p1  *)
          unfold admissible in A3. destruct A3 as [H7 H8]. 

          (* It follows that g u = u *)
          assert (g u = u) as A4. { apply H8, H6. }

          (* It follows that y = u  *)
          assert (y = u) as A5. { rewrite <- A4. symmetry. apply H5. }

          (* So y is free in p1 *)
          assert (y :: Fr p1) as A6. { rewrite A5. apply H6. }

          (* So y is free in All x p1 *)
          assert (y :: Fr (All x p1)) as A7.
          { simpl. apply remove_charac. split.

            - assert (y :: Fr p1) as A. 2:apply A. apply A6.

            - assert (x <> y) as A. 2:apply A. apply not_eq_sym, H4.             
          }
         
          (* Hence from H3 we have f y = y *)
          assert (f y = y) as A8. { apply H3, A7. }

          (* Given that f y = y and y = f x ... *)
          rewrite <- A8, <- E1. apply not_eq_sym.

          (* We therefore need to show that y <> f y ... *) 
          assert (y <> f y) as A. 2: apply A.

          (* ... which follows from H2 ... *)
          apply H2. 

          (* ... provided we show that y is free in All x p1 ...  *)
          assert (y :: Fr (All x p1)) as A. 2: apply A.

          (* ... which has already been  established  *)
          apply A7.

        (* Completes the proof that y is not free in q1 *) 
        } 
Qed.

(* This is a relation which is larger than Alpha0 but a lot simpler. As we      *)
(* shall see, it is also a generator of the alpha-equivalence congruence.       *)
Inductive Alpha1 (v:Type) (e:Eq v) : P v -> P v -> Prop :=
| mkAlpha1: forall (p:P v) (f:v -> v), admissible f p -> Alpha1 v e p (fmap f p)
.

Arguments Alpha1 {v} {e}.
Arguments mkAlpha1 {v} {e}.

(* Alpha-equivalence is also the congruence generated by Alpha1.                *)
Lemma Alpha_admissible_gen : forall (v:Type) (e:Eq v), Alpha = Cong Alpha1.
Proof.
  (* Let v be a Type with decidable equality e  *)
  intros v e.
  
  (* Define r  *)
  remember (Cong Alpha1) as r eqn:E1.

  (* We need to show that Alpha = r *)
  assert (Alpha = r) as A. 2: apply A.

  (* We do so with a double inclusion argument *)
  apply incl_anti.

  (* First we show that Alpha <= r  *)
  - assert (Alpha <= r) as A. 2: apply A.

    (* We argue that Alpha is the smallest congruence containing Alpha0 *)
    unfold Alpha. apply Cong_smallest.

    (* So we need to show that r is a congruence  *)
    + assert (congruence r) as A. 2: apply A.
        
      rewrite E1. apply Cong_congruence.

    (* And we need to show that r contains Alpha0 *)
    + assert (Alpha0 <= r) as A. 2: apply A.

      (* So let x y and p1 such that x <> y and ~ y :: Fr p1  *)
      apply incl_charac. intros p q H1. destruct H1 as [x y p1 H1 H2].

      (* Define p *)
      remember (All x p1) as p eqn:E2.

      (* Define q *)
      remember (All y (fmap (y <:> x) p1)) as q eqn:E3.

      (* Define f *)
      remember (y <:> x) as f eqn:E4.

      (* We need to show that (p,q) :: r  *)
      assert (r p q) as A. 2: apply A.

      (* i.e. that (p.q) belongs to the congruence generated by Alpha1  *)
      rewrite E1. 
        
      (* We argue that (p,q) actually belongs to the generator itself *)
      constructor.

      (* So we need to show that (p,q) belongs to Alpha1  *)
      assert (Alpha1 p q) as A. 2: apply A.

      (* However, q is in fact q = fmap f p *)
      assert (q = fmap f p) as A.
      { rewrite E2, E3. simpl.
        assert (f x = y) as A5. 2: rewrite A5; reflexivity.
        rewrite E4. apply permute_app_right.
      }

      (* So we need to show that (p, fmap f p) lies in Alpha1 *)
      rewrite A. clear A. 
          
      (* which is true by definition... *)
      constructor.  
    
      (* ... provided we show that f is admissible for p  *)
      assert (admissible f p) as A. 2: apply A.
       
      (* Given the definition of an admissible substitution *)
      unfold admissible. split. 

      (* First we need to show that f is valid for p *)
      * assert (valid f p) as A. 2: apply A.
            
        (* It is sufficient to show that f is injective on (var p) *)
        apply valid_inj.
            
        (* It is sufficient to show that f is injective *)
        apply injective_injective_on.

        (* So we now prove that f is injective *)
        assert (injective f) as A. 2: apply A. 
            
        (* However, f is the permutation mapping (y <:> x)  *) 
        rewrite E4. 
            
        (* it is therefore injective  *)
        apply permute_injective.
         

      (* And furthermore that free variables are invariant by f *)
      * assert (forall (u:v), u :: Fr p -> f u = u) as A. 2: apply A.
            
        (* So let u with u :: Fr p  *) 
        intros u H3.
            
        (* We need to show that f u = u *)
        assert (f u = u) as A. 2: apply A.

        (* Given that f is the permutation mapping (y <:> x) ...  *)
        rewrite E4.

        (* ... it is sufficient to show that u <> x and u <> y *)
        apply permute_app_diff. 

        (* First we show that u <> y  *)
        { assert (u <> y) as A. 2: apply A.

          (* Since u :: Fr p, we have u :: Fr p1  *)
          assert (u :: Fr p1) as A.
          { rewrite E2 in H3. simpl in H3.
            apply remove_charac in H3.
            destruct H3 as [H3 H4]. assumption. 
          }
                
          (* So if we assume that u = y ... *)
          intros H4. 

          (* ... we obtain y :: Fr p1 which is a contradiction  *)
          rewrite H4 in A. contradiction. 
        }

        (* We now show that u <> x  *)
        { assert (u <> x) as A. 2: apply A.

          (* This is the case since u is free in p = All x p1 *)
          rewrite E2 in H3. simpl in H3. 
          apply remove_charac in H3.
          destruct H3 as [H3 H4]. apply not_eq_sym.
          assumption.

        } 
          
  (* We now show that r <= Alpha  *)
  - assert (r <= Alpha) as A. 2: apply A.
    
    (* We argue that r is the smallest congruence containing Alpha1 *)
    rewrite E1. apply Cong_smallest.

    (* So we need to show that Alpha is a congruence  *)
    + assert (congruence Alpha) as A. 2: apply A.
      
      unfold Alpha. apply Cong_congruence.
 
    (* And we need to show that Alpha contains Alpha1 *)
    + assert (Alpha1 <= Alpha) as A. 2: apply A.
      
      (* So let p and f : v -> v such that f is admissible for p  *) 
      apply incl_charac. intros p q H5. destruct H5 as [p f H5].

      (* We need to show that p is alpha-equivalent to fmap f p  *)
      assert (p ~ fmap f p) as A. 2: apply A. 

      (* This is the case, provided f is admissible ... *)
      apply Alpha_admissible. 
      
      (* ... which is true by assumption *)
      apply H5. 
Qed.

(* Two alpha-equivalent formulas have the same free variables.                  *)
Lemma Alpha_free : forall (v:Type) (e:Eq v) (p q:P v), 
    p ~ q -> Fr p = Fr q.
Proof.
  (* Let v be a Type with decidable equality e  *)
  intros v e.  

  (* Define r to be the relation 'Fr p = Fr q' *)
  remember (fun (p q:P v) => Fr p = Fr q) as r eqn:E1.

  apply incl_charac. rewrite <- E1.

  (* We need to show that Alpha <= r  *)
  assert (Alpha <= r) as A. 2: apply A.

  (* We argue that Alpha is the smallest congruence containing Alpha1 *)
  rewrite Alpha_admissible_gen. apply Cong_smallest.

  (* So we need to show that r is a congruence ... *)
  - assert (congruence r) as A. 2: apply A.

    rewrite E1. apply free_congruence.

  (* ... and we need to show that r contains Alpha1 *)
  - assert (Alpha1 <= r) as A. 2: apply A.

    (* So let p be a formula and f:v -> v admissible for p *)
    apply incl_charac. intros p q H1. destruct H1 as [p f H1].
    
    (* We need to show that (p, fmap f p) lies in r *)
    assert (r p (fmap f p)) as A. 2: apply A.

    (* Given the way we have defined r ...  *)
    rewrite E1.

    (* ,,, we need to show that p and fmap f p have the same free variables *)
    assert (Fr p = Fr (fmap f p)) as A. 2: apply A.

    (* By transitivity ...  *)
    apply eq_trans with (map f (Fr p)).

    (* ... it is sufiicient to show firstly that Fr p = map f (Fr p) *)
    + assert (Fr p = map f (Fr p)) as A. 2: apply A.

      (* Again by transitivity ... *)
      apply eq_trans with (map id (Fr p)).

      (* ... it is sufficient to show firstly that Fr p = map id (Fr p) *)
      * assert (Fr p = map id (Fr p)) as A. 2: apply A.

        symmetry. apply map_id.

      (* ... and secondly that map id (Fr p) = map f (Fr p) ... *)
      * assert (map id (Fr p) = map f (Fr p)) as A. 2: apply A.

        (* ... which is the case ... *)
        apply coincide_map.

        (* ... provided we show that id and f coincide on Fr p  *)
        assert (coincide (Fr p) id f) as A. 2: apply A.

        (* So let u be a free variable of p *)
        intros u H2.

        (* We need to show that id u = f u *)
        assert (id u = f u) as A. 2: apply A.

        destruct H1 as [H1 H3]. symmetry. apply H3, H2.

    + assert (map f (Fr p) = Fr (fmap f p)) as A. 2: apply A.

      symmetry. destruct H1 as [H1 H3]. 

      apply (valid_free v v e e f p).
        { apply H1. }
        { apply Sub_refl. }
Qed.


(* The binding variable does not matter when not free *) 
Lemma Alpha_not_free_bind : forall (v:Type) (e:Eq v) (p1:P v) (x y:v),
  ~ x :: Fr p1 -> ~ y :: Fr p1 -> All x p1 ~ All y p1. 
Proof.
  (* Let v be a Type with decidable equality e *)
  intros v e.

  (* Let p1 be a formula and x y be variables *)
  intros p1 x y.

  (* We assume that x and y are not free variables of p1 *)
  intros Hx Hy.

  (* We need to distinguish two cases *)
  destruct (eqDec x y) as [H1|H1].

  (* First we assume that x = y *)
  - rewrite <- H1.

    (* We need to show that All x p1 ~ All x p1 *)
    assert (All x p1 ~ All x p1) as A. 2: apply A.

    (* which is true by reflexivity *)
    apply Cong_reflexive.
  
  (* Next we assume that x <> y *)
  -
    (* We need to show that All x p1 is alpha-equivalent to All y p1 *)
    assert (All x p1 ~ All y p1) as A. 2: apply A.

    (* By transitivity, it is sufficient to prove two equivalences *)
    apply Cong_transitive with (All y (fmap (y <:> x) p1)).

    (* First we need to show that All x p1 ~ All y (fmap (y <:> x) p1) *)
    + assert (All x p1 ~ All y (fmap (y <:> x) p1)) as A. 2: apply A.

      (* This is true by definition of alpha-equivalence *)
      constructor. constructor.

      (* since  we have x <> y *)
      * assert (x <> y) as A. 2: apply A. apply H1.

      (* and y is not free in p1 *)
      * assert (~ y :: Fr p1) as A. 2: apply A. apply Hy.

    (* Second we need to show that All y (fmap (y <:> x) p1) ~ All y p1 *)
    + assert (All y (fmap (y <:> x) p1) ~ All y p1) as A. 2: apply A.

      apply CongAll. apply Cong_symmetric.

      (* So it is sufficient to show that fmap (y <:> x) p1 ~ p1 *)
      assert (p1 ~ fmap (y <:> x) p1) as A. 2: apply A.
  
      (* Using lemma Alpha_admissible, it is sufficient to show *)
      apply Alpha_admissible.

      (* that (y <:> x) is admissible for p1 *) 
      assert (admissible (y <:> x) p1) as A. 2: apply A.

      (* which follows from lemma admissible_permute *)
      apply admissible_permute.

        (* and the hypothesis of x y not free in p1 *)
        * assert (~ x :: Fr p1) as A. 2: apply A. apply Hx. 
        * assert (~ y :: Fr p1) as A. 2: apply A. apply Hy.
Qed.

(* Alpha-equivalence is preserved by injective maps *)
Lemma Alpha_injective :
  forall (v w:Type) (e:Eq v) (e':Eq w) (f:v -> w) (p q:P v),
    injective f -> p ~ q -> fmap f p ~ fmap f q.
Proof.
  (* Let v w be types with respective decidable equality e e' *)
  intros v w e e'.

  (* Let f be a map from v to w and p q be formulas *)
  intros f p q.

  (* We assume that f is injective *)
  intros HInj. assert (injective f) as A. apply HInj. clear A.

  (* We need to show the implication p ~ q -> fmap f p ~ fmap f q *)
  assert (p ~ q -> fmap f p ~ fmap f q) as A. 2: apply A.

  (* Define the relation r as r p q = fmap f p ~ fmap f q *)
  remember (fun (p q:P v) => fmap f p ~ fmap f q) as r eqn:Er.

  (* Then r p q = fmap f p ~ fmap f q *)
  assert (r p q = fmap f p ~ fmap f q) as E. rewrite Er. reflexivity.

  (* So we need to show the implication p ~ q -> r p q for all p q *)
  rewrite <- E. clear E. revert q. revert p.
  assert (forall (p q:P v), p ~ q -> r p q) as A. 2: apply A.

  (* In other words, we need to show thw inclusion ~ <= r *)
  rewrite <- incl_charac.
  assert (Alpha <= r) as A. 2: apply A.

  (* Alpha being the smallest congruence on P v which contains Alpha0 *)
  apply Cong_smallest.

  (* It is sufficient first show that r is a congruence on P v *)
  - assert (congruence r) as A. 2: apply A. 

    (* which follows from Lemma fmap_congruence *)
    rewrite Er. apply fmap_congruence.

    (* together with the fact that alpha-equivalence is itself a congruence *)
    assert (congruence Alpha) as A. 2: apply A.

    (* which is true since Alpha is the congruence generated by Alpha0 *)
    apply Cong_congruence.

  (* and second to show that r contains Alpha0 *)
  - assert (Alpha0 <= r) as A. 2: apply A.

    (* So let x y be variables and p1 be a formula *)
    rewrite incl_charac.
    intros p' q' H. destruct H as [x y p1 H3 H4]. 

    (* such that x <> y *)
    assert (x <> y) as A. apply H3. clear A. 

    (* and y is not free in p1 *)
    assert (~ y :: Fr p1) as A. apply H4. clear A.

    (* Define p = All x p1 *)
    remember (All x p1) as p eqn:Ep.

    (* Define q = All y (fmap (y <:> x) p1) *)
    remember (All y (fmap (y <:> x) p1)) as q eqn:Eq.

    (* Then we simply need to show that r p q holds *)
    assert (r p q) as A. 2: apply A.

    (* or in other words that fmap f p ~ fmap f q *)
    rewrite Er.
    assert (fmap f p ~ fmap f q) as A. 2: apply A.

    (* It is sufficient to show that Alpha0 (fmap f p) (fmap f q) *)
    apply CongBase.
    assert (Alpha0 (fmap f p) (fmap f q)) as A. 2: apply A.

    (* So it is sufficient to show the existence of p1' : P w
       and x' y' : w with x' <> y' and y' not free in p1' such that
       fmap f p = All x' p1' and fmap f q = All y' (fmap (y'<:>x') p1') *)
    
    (* Define p1' = fmap f p1 *)
    remember (fmap f p1) as p1' eqn:Ep1'.
    
    (* Define x' = f x *)
    remember (f x) as x' eqn:Ex'.

    (* Define y' = f y *)
    remember (f y) as y' eqn:Ey'.

    (* Then we do have fmap f p = All x' p1' *)
    assert (fmap f p = All x' p1') as E1.
      { rewrite Ep, Ex', Ep1'. reflexivity. }

    (* and fmap f q = All y' (fmap <y':x'> p1') *)
    assert (fmap f q = All y' (fmap (y'<:>x') p1')) as E2.
      { rewrite Eq, Ex', Ey', Ep1'. simpl.
        rewrite <- fmap_comp', <- fmap_comp'.
        rewrite <- (permute_comp v w e e'). 
        reflexivity. 
        apply HInj. (* f is injective *)
      }

    (* we also have x' <> y' *)
    assert (x' <> y') as HNeq.
      { rewrite Ex', Ey'. intro H. apply HInj in H. contradiction. } 

    (* and y' is not free in p1' *)
    assert (~ y' :: Fr p1') as HFree.
    { rewrite Ep1'. rewrite (free_inj v w e e'). 
      2: apply injective_injective_on, HInj.
      intro HFree. apply in_map_iff in HFree. 
      destruct HFree as [u [H1 H2]].
      rewrite Ey' in H1. apply HInj in H1. subst. 
      contradiction.
    }

    (* which allows us to conclude *)
    rewrite E1,E2. constructor.
      { apply HNeq. }
      { apply HFree. }
Qed.
