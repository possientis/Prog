Require Import List.

Require Import Logic.Class.Eq.

Require Import Logic.Func.Permute.
Require Import Logic.Func.Identity.
Require Import Logic.Func.Injective.
Require Import Logic.Func.Composition.

Require Import Logic.List.In.
Require Import Logic.List.Remove.
Require Import Logic.List.Append.
Require Import Logic.List.InjectiveOn.

Require Import Logic.Fol.Free.
Require Import Logic.Fol.Valid.
Require Import Logic.Fol.Syntax.
Require Import Logic.Fol.Functor.
Require Import Logic.Fol.Variable.
Require Import Logic.Fol.Congruence.
Require Import Logic.Fol.Admissible.

(* Generator of alpha-equivalence.                                              *)
(* We wish to formally define alpha-equivalence as the smallest congruence      *)
(* contaning all ordered pairs below. Note that we are using the permutation    *)
(* y <:> x rather than the substitution (y // x) and we allow the variable y    *)
(* to be a variable of p1 as long as it is not free. This seemingly unusual     *)
(* choice is to make sure we obtain a definition of alpha-equivalence which     *)
(* works equally well for a finite or infinite variable type v. Otherwise, we   *)
(* would obtain a congruence which is strictly stronger than alpha-equivalence  *)
(* when v is finite. See the StrongAlpha module for details.                    *)
Inductive Alpha0 (v:Type) (e:Eq v) : P v -> P v -> Prop :=
| mkAlpha0: forall (x y:v) (p1:P v), 
    x <> y       -> 
    ~ y :: Fr p1 ->
    Alpha0 v e (All x p1) (All y (fmap (y <:> x) p1)) 
.

Arguments Alpha0 {v} {e}.
Arguments mkAlpha0 {v} {e}.

(* The alpha-equivalence relation is the congruence generated by Alph0.         *)
Definition Alpha (v:Type) (e:Eq v) : P v -> P v -> Prop := 
    Cong (@Alpha0 v e).

Arguments Alpha {v} {e}.

Notation "p ~ q" := (Alpha p q)
    (at level 60, no associativity) : Fol_Alpha_scope.

Open Scope Fol_Alpha_scope.

(* Admissible substitutions do not change alpha-equivalence classes.            *)
Lemma Alpha_admissible : forall (v:Type) (e:Eq v) (p:P v) (f:v -> v),
  admissible f p -> p ~ fmap f p.
Proof.
  intros v e.
  induction p as [|x y|p1 IH1 p2 IH2|x p1 IH1]; 
  intros f [H1 H2]; simpl; simpl in H2.

  (* case p = Bot *)
  - apply Cong_reflexive.

  (* case p = Elem x y *)
  - assert (f x = x) as E1. { apply H2. left. reflexivity. }
    assert (f y = y) as E2. { apply H2. right. left. reflexivity. }
    rewrite E1, E2. apply Cong_reflexive.

  (* case p = Imp p1 p2 *)
  - rewrite valid_imp in H1; destruct H1 as [H1 H3].

    assert (p1 ~ fmap f p1) as E1.
      { apply IH1. unfold admissible. split.
        { assumption. }
        { intros x H4. apply H2, app_charac. left. assumption. }}

    assert (p2 ~ fmap f p2) as E2.
      { apply IH2. unfold admissible. split.
        { assumption. }
        { intros x H4. apply H2, app_charac. right. assumption. }}

    apply CongImp; assumption. 

  (* case p = All x p1 *)
  - rewrite valid_all in H1. destruct H1 as [H3 H4].
    destruct (eqDec (f x) x) as [H5|H5].

    + (* f x = x *)
      assert (p1 ~ fmap f p1) as E1.
        { apply IH1. unfold admissible. split.
          { assumption. }
          { intros y H6.
            assert (f y = y) as E1.
              { destruct (eqDec x y) as [H7|H7].
                { (* x = y  *)
                  rewrite <- H7. assumption. }
                { (* x <> y *)
                  apply H2, remove_charac. split; assumption. }}
           assumption. }} 
      rewrite H5. apply CongAll. assumption.

    + (* f x <> x *)
      remember (f x) as y eqn:H6.

      assert (All x p1 ~ All y (fmap f p1)) as E.
        { remember ((y <:> x) ; f) as g eqn:H7.
          remember (fmap g p1) as q1 eqn:H8. 

          assert (f = (y <:> x) ; g) as E1.
            { rewrite H7. rewrite comp_assoc, permute_involution.
              symmetry. apply comp_id_left. }

          assert (fmap f p1 = fmap (y <:> x) q1) as E2.
            { rewrite H8, <- fmap_comp', <- E1. reflexivity. }

          rewrite E2.

          assert (All x p1 ~ All y (fmap (y <:> x) q1)) as E3.
            { assert (admissible g p1) as E8. 
                { unfold admissible. split.
                  { rewrite H7. rewrite <- valid_compose. split.
                    { apply H3. (* why is the assumption tactic failing here *) }
                    { apply valid_inj, injective_injective_on. 
                      apply permute_injective. }}
                  { intros u H10. destruct (eqDec u x) as [H11|H11].
                    { subst. unfold comp. apply permute_app_left. }
                    { rewrite H7. unfold comp. 
                      assert (f u = u) as H12.
                        { apply H2. apply remove_charac. split.
                          { assumption. }
                          { intros H12. apply H11. symmetry.  assumption. }}
                      rewrite H12. apply permute_app_diff. 
                        { intros H13. apply H4 with u. 
                          { simpl. apply remove_charac. split.
                            { assumption. }
                            { intros H14. apply H11. symmetry. assumption. }}
                          { rewrite H12. symmetry. assumption. }}
                        { assumption. }}}}

              assert (~ y :: Fr q1) as E4.
                { rewrite H8. intros H9. apply (free_fmap v v e) in H9.
                  apply in_map_iff in H9. destruct H9 as [u [H9 H10]].
                  unfold admissible in E8. destruct E8 as [H11 H12]. 

                  assert (g u = u) as H13. { apply H12. assumption. }

                  assert (y :: Fr p1) as H14. { rewrite <- H9, H13. assumption. }

                  assert (y :: Fr (All x p1)) as H15.
                    { simpl. apply remove_charac. split.
                      { assumption. }
                      { intros H16. apply H5. symmetry. assumption. }} 

                  assert (f y = y) as H17. { apply H2. assumption. }

                  assert (f x <> f y) as H18. 
                    { rewrite <- H6. apply H4. assumption. }

                  assert (f x <> y) as H19. { rewrite <- H17. assumption. }

                  apply H19. symmetry. assumption. }

              assert (All x q1 ~ All y (fmap (y <:> x) q1)) as E5.
                { constructor. constructor.
                  { intros H9. apply H5. symmetry. assumption. }
                  { assumption. }}

              assert (All x p1 ~ All x q1) as E6.
                { assert (p1 ~ q1) as E7. { rewrite H8. apply IH1. apply E8. }
                  apply Cong_congruent, E7. }

              apply Cong_transitive with (All x q1); assumption. }
          apply E3. }
      apply E.
Qed.

